VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_2_16_sky130A
   CLASS BLOCK ;
   SIZE 108.31 BY 121.23 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  10.69 -10.39 11.07 -10.01 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  22.25 -10.39 22.63 -10.01 ;
      END
   END din0[1]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -11.75 120.85 -11.37 121.23 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -13.79 120.85 -13.41 121.23 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -12.43 120.85 -12.05 121.23 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -13.11 120.85 -12.73 121.23 ;
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  -104.23 -7.67 -103.85 -7.29 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  -104.23 -3.59 -103.85 -3.21 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -57.99 -10.39 -57.61 -10.01 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m3 ;
         RECT  107.93 11.37 108.31 11.75 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m3 ;
         RECT  107.93 10.01 108.31 10.39 ;
      END
   END dout0[1]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  -103.55 -5.63 -102.49 -4.57 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  -104.23 -9.71 -103.17 -9.33 ;
      END
   END gnd
   OBS
   LAYER  m1 ;
      RECT  92.53 37.14 92.82 37.43 ;
      RECT  92.98 34.54 93.3 34.86 ;
      RECT  91.79 35.02 92.12 35.17 ;
      RECT  92.47 34.54 92.79 34.86 ;
      RECT  92.95 37.68 93.24 37.97 ;
      RECT  91.61 39.04 94.21 39.33 ;
      RECT  91.81 35.17 92.1 35.33 ;
      RECT  91.61 33.96 94.21 34.25 ;
      RECT  92.53 41.24 92.82 40.95 ;
      RECT  92.98 43.84 93.3 43.52 ;
      RECT  91.79 43.36 92.12 43.21 ;
      RECT  92.47 43.84 92.79 43.52 ;
      RECT  92.95 40.7 93.24 40.41 ;
      RECT  91.61 39.34 94.21 39.05 ;
      RECT  91.81 43.21 92.1 43.05 ;
      RECT  91.61 44.42 94.21 44.13 ;
      RECT  92.53 47.32 92.82 47.61 ;
      RECT  92.98 44.72 93.3 45.04 ;
      RECT  91.79 45.2 92.12 45.35 ;
      RECT  92.47 44.72 92.79 45.04 ;
      RECT  92.95 47.86 93.24 48.15 ;
      RECT  91.61 49.22 94.21 49.51 ;
      RECT  91.81 45.35 92.1 45.51 ;
      RECT  91.61 44.14 94.21 44.43 ;
      RECT  92.53 51.42 92.82 51.13 ;
      RECT  92.98 54.02 93.3 53.7 ;
      RECT  91.79 53.54 92.12 53.39 ;
      RECT  92.47 54.02 92.79 53.7 ;
      RECT  92.95 50.88 93.24 50.59 ;
      RECT  91.61 49.52 94.21 49.23 ;
      RECT  91.81 53.39 92.1 53.23 ;
      RECT  91.61 54.6 94.21 54.31 ;
      RECT  92.53 57.5 92.82 57.79 ;
      RECT  92.98 54.9 93.3 55.22 ;
      RECT  91.79 55.38 92.12 55.53 ;
      RECT  92.47 54.9 92.79 55.22 ;
      RECT  92.95 58.04 93.24 58.33 ;
      RECT  91.61 59.4 94.21 59.69 ;
      RECT  91.81 55.53 92.1 55.69 ;
      RECT  91.61 54.32 94.21 54.61 ;
      RECT  92.53 61.6 92.82 61.31 ;
      RECT  92.98 64.2 93.3 63.88 ;
      RECT  91.79 63.72 92.12 63.57 ;
      RECT  92.47 64.2 92.79 63.88 ;
      RECT  92.95 61.06 93.24 60.77 ;
      RECT  91.61 59.7 94.21 59.41 ;
      RECT  91.81 63.57 92.1 63.41 ;
      RECT  91.61 64.78 94.21 64.49 ;
      RECT  92.53 67.68 92.82 67.97 ;
      RECT  92.98 65.08 93.3 65.4 ;
      RECT  91.79 65.56 92.12 65.71 ;
      RECT  92.47 65.08 92.79 65.4 ;
      RECT  92.95 68.22 93.24 68.51 ;
      RECT  91.61 69.58 94.21 69.87 ;
      RECT  91.81 65.71 92.1 65.87 ;
      RECT  91.61 64.5 94.21 64.79 ;
      RECT  92.53 71.78 92.82 71.49 ;
      RECT  92.98 74.38 93.3 74.06 ;
      RECT  91.79 73.9 92.12 73.75 ;
      RECT  92.47 74.38 92.79 74.06 ;
      RECT  92.95 71.24 93.24 70.95 ;
      RECT  91.61 69.88 94.21 69.59 ;
      RECT  91.81 73.75 92.1 73.59 ;
      RECT  91.61 74.96 94.21 74.67 ;
      RECT  92.53 77.86 92.82 78.15 ;
      RECT  92.98 75.26 93.3 75.58 ;
      RECT  91.79 75.74 92.12 75.89 ;
      RECT  92.47 75.26 92.79 75.58 ;
      RECT  92.95 78.4 93.24 78.69 ;
      RECT  91.61 79.76 94.21 80.05 ;
      RECT  91.81 75.89 92.1 76.05 ;
      RECT  91.61 74.68 94.21 74.97 ;
      RECT  92.53 81.96 92.82 81.67 ;
      RECT  92.98 84.56 93.3 84.24 ;
      RECT  91.79 84.08 92.12 83.93 ;
      RECT  92.47 84.56 92.79 84.24 ;
      RECT  92.95 81.42 93.24 81.13 ;
      RECT  91.61 80.06 94.21 79.77 ;
      RECT  91.81 83.93 92.1 83.77 ;
      RECT  91.61 85.14 94.21 84.85 ;
      RECT  92.53 88.04 92.82 88.33 ;
      RECT  92.98 85.44 93.3 85.76 ;
      RECT  91.79 85.92 92.12 86.07 ;
      RECT  92.47 85.44 92.79 85.76 ;
      RECT  92.95 88.58 93.24 88.87 ;
      RECT  91.61 89.94 94.21 90.23 ;
      RECT  91.81 86.07 92.1 86.23 ;
      RECT  91.61 84.86 94.21 85.15 ;
      RECT  92.53 92.14 92.82 91.85 ;
      RECT  92.98 94.74 93.3 94.42 ;
      RECT  91.79 94.26 92.12 94.11 ;
      RECT  92.47 94.74 92.79 94.42 ;
      RECT  92.95 91.6 93.24 91.31 ;
      RECT  91.61 90.24 94.21 89.95 ;
      RECT  91.81 94.11 92.1 93.95 ;
      RECT  91.61 95.32 94.21 95.03 ;
      RECT  92.53 98.22 92.82 98.51 ;
      RECT  92.98 95.62 93.3 95.94 ;
      RECT  91.79 96.1 92.12 96.25 ;
      RECT  92.47 95.62 92.79 95.94 ;
      RECT  92.95 98.76 93.24 99.05 ;
      RECT  91.61 100.12 94.21 100.41 ;
      RECT  91.81 96.25 92.1 96.41 ;
      RECT  91.61 95.04 94.21 95.33 ;
      RECT  92.53 102.32 92.82 102.03 ;
      RECT  92.98 104.92 93.3 104.6 ;
      RECT  91.79 104.44 92.12 104.29 ;
      RECT  92.47 104.92 92.79 104.6 ;
      RECT  92.95 101.78 93.24 101.49 ;
      RECT  91.61 100.42 94.21 100.13 ;
      RECT  91.81 104.29 92.1 104.13 ;
      RECT  91.61 105.5 94.21 105.21 ;
      RECT  92.53 108.4 92.82 108.69 ;
      RECT  92.98 105.8 93.3 106.12 ;
      RECT  91.79 106.28 92.12 106.43 ;
      RECT  92.47 105.8 92.79 106.12 ;
      RECT  92.95 108.94 93.24 109.23 ;
      RECT  91.61 110.3 94.21 110.59 ;
      RECT  91.81 106.43 92.1 106.59 ;
      RECT  91.61 105.22 94.21 105.51 ;
      RECT  92.53 112.5 92.82 112.21 ;
      RECT  92.98 115.1 93.3 114.78 ;
      RECT  91.79 114.62 92.12 114.47 ;
      RECT  92.47 115.1 92.79 114.78 ;
      RECT  92.95 111.96 93.24 111.67 ;
      RECT  91.61 110.6 94.21 110.31 ;
      RECT  91.81 114.47 92.1 114.31 ;
      RECT  91.61 115.68 94.21 115.39 ;
      RECT  95.13 37.14 95.42 37.43 ;
      RECT  95.58 34.54 95.9 34.86 ;
      RECT  94.39 35.02 94.72 35.17 ;
      RECT  95.07 34.54 95.39 34.86 ;
      RECT  95.55 37.68 95.84 37.97 ;
      RECT  94.21 39.04 96.81 39.33 ;
      RECT  94.41 35.17 94.7 35.33 ;
      RECT  94.21 33.96 96.81 34.25 ;
      RECT  95.13 41.24 95.42 40.95 ;
      RECT  95.58 43.84 95.9 43.52 ;
      RECT  94.39 43.36 94.72 43.21 ;
      RECT  95.07 43.84 95.39 43.52 ;
      RECT  95.55 40.7 95.84 40.41 ;
      RECT  94.21 39.34 96.81 39.05 ;
      RECT  94.41 43.21 94.7 43.05 ;
      RECT  94.21 44.42 96.81 44.13 ;
      RECT  95.13 47.32 95.42 47.61 ;
      RECT  95.58 44.72 95.9 45.04 ;
      RECT  94.39 45.2 94.72 45.35 ;
      RECT  95.07 44.72 95.39 45.04 ;
      RECT  95.55 47.86 95.84 48.15 ;
      RECT  94.21 49.22 96.81 49.51 ;
      RECT  94.41 45.35 94.7 45.51 ;
      RECT  94.21 44.14 96.81 44.43 ;
      RECT  95.13 51.42 95.42 51.13 ;
      RECT  95.58 54.02 95.9 53.7 ;
      RECT  94.39 53.54 94.72 53.39 ;
      RECT  95.07 54.02 95.39 53.7 ;
      RECT  95.55 50.88 95.84 50.59 ;
      RECT  94.21 49.52 96.81 49.23 ;
      RECT  94.41 53.39 94.7 53.23 ;
      RECT  94.21 54.6 96.81 54.31 ;
      RECT  95.13 57.5 95.42 57.79 ;
      RECT  95.58 54.9 95.9 55.22 ;
      RECT  94.39 55.38 94.72 55.53 ;
      RECT  95.07 54.9 95.39 55.22 ;
      RECT  95.55 58.04 95.84 58.33 ;
      RECT  94.21 59.4 96.81 59.69 ;
      RECT  94.41 55.53 94.7 55.69 ;
      RECT  94.21 54.32 96.81 54.61 ;
      RECT  95.13 61.6 95.42 61.31 ;
      RECT  95.58 64.2 95.9 63.88 ;
      RECT  94.39 63.72 94.72 63.57 ;
      RECT  95.07 64.2 95.39 63.88 ;
      RECT  95.55 61.06 95.84 60.77 ;
      RECT  94.21 59.7 96.81 59.41 ;
      RECT  94.41 63.57 94.7 63.41 ;
      RECT  94.21 64.78 96.81 64.49 ;
      RECT  95.13 67.68 95.42 67.97 ;
      RECT  95.58 65.08 95.9 65.4 ;
      RECT  94.39 65.56 94.72 65.71 ;
      RECT  95.07 65.08 95.39 65.4 ;
      RECT  95.55 68.22 95.84 68.51 ;
      RECT  94.21 69.58 96.81 69.87 ;
      RECT  94.41 65.71 94.7 65.87 ;
      RECT  94.21 64.5 96.81 64.79 ;
      RECT  95.13 71.78 95.42 71.49 ;
      RECT  95.58 74.38 95.9 74.06 ;
      RECT  94.39 73.9 94.72 73.75 ;
      RECT  95.07 74.38 95.39 74.06 ;
      RECT  95.55 71.24 95.84 70.95 ;
      RECT  94.21 69.88 96.81 69.59 ;
      RECT  94.41 73.75 94.7 73.59 ;
      RECT  94.21 74.96 96.81 74.67 ;
      RECT  95.13 77.86 95.42 78.15 ;
      RECT  95.58 75.26 95.9 75.58 ;
      RECT  94.39 75.74 94.72 75.89 ;
      RECT  95.07 75.26 95.39 75.58 ;
      RECT  95.55 78.4 95.84 78.69 ;
      RECT  94.21 79.76 96.81 80.05 ;
      RECT  94.41 75.89 94.7 76.05 ;
      RECT  94.21 74.68 96.81 74.97 ;
      RECT  95.13 81.96 95.42 81.67 ;
      RECT  95.58 84.56 95.9 84.24 ;
      RECT  94.39 84.08 94.72 83.93 ;
      RECT  95.07 84.56 95.39 84.24 ;
      RECT  95.55 81.42 95.84 81.13 ;
      RECT  94.21 80.06 96.81 79.77 ;
      RECT  94.41 83.93 94.7 83.77 ;
      RECT  94.21 85.14 96.81 84.85 ;
      RECT  95.13 88.04 95.42 88.33 ;
      RECT  95.58 85.44 95.9 85.76 ;
      RECT  94.39 85.92 94.72 86.07 ;
      RECT  95.07 85.44 95.39 85.76 ;
      RECT  95.55 88.58 95.84 88.87 ;
      RECT  94.21 89.94 96.81 90.23 ;
      RECT  94.41 86.07 94.7 86.23 ;
      RECT  94.21 84.86 96.81 85.15 ;
      RECT  95.13 92.14 95.42 91.85 ;
      RECT  95.58 94.74 95.9 94.42 ;
      RECT  94.39 94.26 94.72 94.11 ;
      RECT  95.07 94.74 95.39 94.42 ;
      RECT  95.55 91.6 95.84 91.31 ;
      RECT  94.21 90.24 96.81 89.95 ;
      RECT  94.41 94.11 94.7 93.95 ;
      RECT  94.21 95.32 96.81 95.03 ;
      RECT  95.13 98.22 95.42 98.51 ;
      RECT  95.58 95.62 95.9 95.94 ;
      RECT  94.39 96.1 94.72 96.25 ;
      RECT  95.07 95.62 95.39 95.94 ;
      RECT  95.55 98.76 95.84 99.05 ;
      RECT  94.21 100.12 96.81 100.41 ;
      RECT  94.41 96.25 94.7 96.41 ;
      RECT  94.21 95.04 96.81 95.33 ;
      RECT  95.13 102.32 95.42 102.03 ;
      RECT  95.58 104.92 95.9 104.6 ;
      RECT  94.39 104.44 94.72 104.29 ;
      RECT  95.07 104.92 95.39 104.6 ;
      RECT  95.55 101.78 95.84 101.49 ;
      RECT  94.21 100.42 96.81 100.13 ;
      RECT  94.41 104.29 94.7 104.13 ;
      RECT  94.21 105.5 96.81 105.21 ;
      RECT  95.13 108.4 95.42 108.69 ;
      RECT  95.58 105.8 95.9 106.12 ;
      RECT  94.39 106.28 94.72 106.43 ;
      RECT  95.07 105.8 95.39 106.12 ;
      RECT  95.55 108.94 95.84 109.23 ;
      RECT  94.21 110.3 96.81 110.59 ;
      RECT  94.41 106.43 94.7 106.59 ;
      RECT  94.21 105.22 96.81 105.51 ;
      RECT  95.13 112.5 95.42 112.21 ;
      RECT  95.58 115.1 95.9 114.78 ;
      RECT  94.39 114.62 94.72 114.47 ;
      RECT  95.07 115.1 95.39 114.78 ;
      RECT  95.55 111.96 95.84 111.67 ;
      RECT  94.21 110.6 96.81 110.31 ;
      RECT  94.41 114.47 94.7 114.31 ;
      RECT  94.21 115.68 96.81 115.39 ;
      RECT  91.61 35.17 96.81 35.33 ;
      RECT  91.61 43.05 96.81 43.21 ;
      RECT  91.61 45.35 96.81 45.51 ;
      RECT  91.61 53.23 96.81 53.39 ;
      RECT  91.61 55.53 96.81 55.69 ;
      RECT  91.61 63.41 96.81 63.57 ;
      RECT  91.61 65.71 96.81 65.87 ;
      RECT  91.61 73.59 96.81 73.75 ;
      RECT  91.61 75.89 96.81 76.05 ;
      RECT  91.61 83.77 96.81 83.93 ;
      RECT  91.61 86.07 96.81 86.23 ;
      RECT  91.61 93.95 96.81 94.11 ;
      RECT  91.61 96.25 96.81 96.41 ;
      RECT  91.61 104.13 96.81 104.29 ;
      RECT  91.61 106.43 96.81 106.59 ;
      RECT  91.61 114.31 96.81 114.47 ;
      RECT  91.61 110.31 94.21 110.6 ;
      RECT  94.21 110.31 96.81 110.6 ;
      RECT  94.21 39.04 96.81 39.33 ;
      RECT  94.21 79.76 96.81 80.05 ;
      RECT  94.21 89.94 96.81 90.23 ;
      RECT  91.61 89.95 94.21 90.24 ;
      RECT  91.61 79.76 94.21 80.05 ;
      RECT  94.21 69.58 96.81 69.87 ;
      RECT  94.21 89.95 96.81 90.24 ;
      RECT  91.61 79.77 94.21 80.06 ;
      RECT  94.21 59.41 96.81 59.7 ;
      RECT  91.61 59.4 94.21 59.69 ;
      RECT  94.21 49.23 96.81 49.52 ;
      RECT  94.21 59.4 96.81 59.69 ;
      RECT  91.61 110.3 94.21 110.59 ;
      RECT  94.21 110.3 96.81 110.59 ;
      RECT  91.61 49.23 94.21 49.52 ;
      RECT  94.21 49.22 96.81 49.51 ;
      RECT  94.21 69.59 96.81 69.88 ;
      RECT  91.61 100.12 94.21 100.41 ;
      RECT  91.61 100.13 94.21 100.42 ;
      RECT  91.61 49.22 94.21 49.51 ;
      RECT  91.61 69.58 94.21 69.87 ;
      RECT  94.21 100.13 96.81 100.42 ;
      RECT  94.21 100.12 96.81 100.41 ;
      RECT  94.21 79.77 96.81 80.06 ;
      RECT  91.61 69.59 94.21 69.88 ;
      RECT  91.61 39.04 94.21 39.33 ;
      RECT  94.21 39.05 96.81 39.34 ;
      RECT  91.61 39.05 94.21 39.34 ;
      RECT  91.61 59.41 94.21 59.7 ;
      RECT  91.61 89.94 94.21 90.23 ;
      RECT  91.61 74.68 94.21 74.97 ;
      RECT  94.21 105.22 96.81 105.51 ;
      RECT  91.61 74.67 94.21 74.96 ;
      RECT  91.61 105.21 94.21 105.5 ;
      RECT  91.61 33.96 94.21 34.25 ;
      RECT  94.21 44.14 96.81 44.43 ;
      RECT  94.21 44.13 96.81 44.42 ;
      RECT  94.21 64.5 96.81 64.79 ;
      RECT  91.61 44.14 94.21 44.43 ;
      RECT  91.61 54.32 94.21 54.61 ;
      RECT  91.61 95.03 94.21 95.32 ;
      RECT  91.61 64.49 94.21 64.78 ;
      RECT  94.21 33.96 96.81 34.25 ;
      RECT  94.21 95.04 96.81 95.33 ;
      RECT  91.61 115.39 94.21 115.68 ;
      RECT  91.61 64.5 94.21 64.79 ;
      RECT  94.21 84.85 96.81 85.14 ;
      RECT  94.21 84.86 96.81 85.15 ;
      RECT  91.61 54.31 94.21 54.6 ;
      RECT  94.21 115.39 96.81 115.68 ;
      RECT  91.61 105.22 94.21 105.51 ;
      RECT  94.21 105.21 96.81 105.5 ;
      RECT  94.21 54.31 96.81 54.6 ;
      RECT  94.21 74.68 96.81 74.97 ;
      RECT  91.61 84.85 94.21 85.14 ;
      RECT  91.61 84.86 94.21 85.15 ;
      RECT  94.21 64.49 96.81 64.78 ;
      RECT  91.61 44.13 94.21 44.42 ;
      RECT  94.21 74.67 96.81 74.96 ;
      RECT  94.21 95.03 96.81 95.32 ;
      RECT  91.61 95.04 94.21 95.33 ;
      RECT  94.21 54.32 96.81 54.61 ;
      RECT  89.93 26.96 90.22 27.25 ;
      RECT  90.38 24.36 90.7 24.68 ;
      RECT  89.19 24.84 89.52 24.99 ;
      RECT  89.87 24.36 90.19 24.68 ;
      RECT  90.35 27.5 90.64 27.79 ;
      RECT  89.01 28.86 91.61 29.15 ;
      RECT  89.21 24.99 89.5 25.15 ;
      RECT  89.01 23.78 91.61 24.07 ;
      RECT  89.93 31.06 90.22 30.77 ;
      RECT  90.38 33.66 90.7 33.34 ;
      RECT  89.19 33.18 89.52 33.03 ;
      RECT  89.87 33.66 90.19 33.34 ;
      RECT  90.35 30.52 90.64 30.23 ;
      RECT  89.01 29.16 91.61 28.87 ;
      RECT  89.21 33.03 89.5 32.87 ;
      RECT  89.01 34.24 91.61 33.95 ;
      RECT  89.93 37.14 90.22 37.43 ;
      RECT  90.38 34.54 90.7 34.86 ;
      RECT  89.19 35.02 89.52 35.17 ;
      RECT  89.87 34.54 90.19 34.86 ;
      RECT  90.35 37.68 90.64 37.97 ;
      RECT  89.01 39.04 91.61 39.33 ;
      RECT  89.21 35.17 89.5 35.33 ;
      RECT  89.01 33.96 91.61 34.25 ;
      RECT  89.93 41.24 90.22 40.95 ;
      RECT  90.38 43.84 90.7 43.52 ;
      RECT  89.19 43.36 89.52 43.21 ;
      RECT  89.87 43.84 90.19 43.52 ;
      RECT  90.35 40.7 90.64 40.41 ;
      RECT  89.01 39.34 91.61 39.05 ;
      RECT  89.21 43.21 89.5 43.05 ;
      RECT  89.01 44.42 91.61 44.13 ;
      RECT  89.93 47.32 90.22 47.61 ;
      RECT  90.38 44.72 90.7 45.04 ;
      RECT  89.19 45.2 89.52 45.35 ;
      RECT  89.87 44.72 90.19 45.04 ;
      RECT  90.35 47.86 90.64 48.15 ;
      RECT  89.01 49.22 91.61 49.51 ;
      RECT  89.21 45.35 89.5 45.51 ;
      RECT  89.01 44.14 91.61 44.43 ;
      RECT  89.93 51.42 90.22 51.13 ;
      RECT  90.38 54.02 90.7 53.7 ;
      RECT  89.19 53.54 89.52 53.39 ;
      RECT  89.87 54.02 90.19 53.7 ;
      RECT  90.35 50.88 90.64 50.59 ;
      RECT  89.01 49.52 91.61 49.23 ;
      RECT  89.21 53.39 89.5 53.23 ;
      RECT  89.01 54.6 91.61 54.31 ;
      RECT  89.93 57.5 90.22 57.79 ;
      RECT  90.38 54.9 90.7 55.22 ;
      RECT  89.19 55.38 89.52 55.53 ;
      RECT  89.87 54.9 90.19 55.22 ;
      RECT  90.35 58.04 90.64 58.33 ;
      RECT  89.01 59.4 91.61 59.69 ;
      RECT  89.21 55.53 89.5 55.69 ;
      RECT  89.01 54.32 91.61 54.61 ;
      RECT  89.93 61.6 90.22 61.31 ;
      RECT  90.38 64.2 90.7 63.88 ;
      RECT  89.19 63.72 89.52 63.57 ;
      RECT  89.87 64.2 90.19 63.88 ;
      RECT  90.35 61.06 90.64 60.77 ;
      RECT  89.01 59.7 91.61 59.41 ;
      RECT  89.21 63.57 89.5 63.41 ;
      RECT  89.01 64.78 91.61 64.49 ;
      RECT  89.93 67.68 90.22 67.97 ;
      RECT  90.38 65.08 90.7 65.4 ;
      RECT  89.19 65.56 89.52 65.71 ;
      RECT  89.87 65.08 90.19 65.4 ;
      RECT  90.35 68.22 90.64 68.51 ;
      RECT  89.01 69.58 91.61 69.87 ;
      RECT  89.21 65.71 89.5 65.87 ;
      RECT  89.01 64.5 91.61 64.79 ;
      RECT  89.93 71.78 90.22 71.49 ;
      RECT  90.38 74.38 90.7 74.06 ;
      RECT  89.19 73.9 89.52 73.75 ;
      RECT  89.87 74.38 90.19 74.06 ;
      RECT  90.35 71.24 90.64 70.95 ;
      RECT  89.01 69.88 91.61 69.59 ;
      RECT  89.21 73.75 89.5 73.59 ;
      RECT  89.01 74.96 91.61 74.67 ;
      RECT  89.93 77.86 90.22 78.15 ;
      RECT  90.38 75.26 90.7 75.58 ;
      RECT  89.19 75.74 89.52 75.89 ;
      RECT  89.87 75.26 90.19 75.58 ;
      RECT  90.35 78.4 90.64 78.69 ;
      RECT  89.01 79.76 91.61 80.05 ;
      RECT  89.21 75.89 89.5 76.05 ;
      RECT  89.01 74.68 91.61 74.97 ;
      RECT  89.93 81.96 90.22 81.67 ;
      RECT  90.38 84.56 90.7 84.24 ;
      RECT  89.19 84.08 89.52 83.93 ;
      RECT  89.87 84.56 90.19 84.24 ;
      RECT  90.35 81.42 90.64 81.13 ;
      RECT  89.01 80.06 91.61 79.77 ;
      RECT  89.21 83.93 89.5 83.77 ;
      RECT  89.01 85.14 91.61 84.85 ;
      RECT  89.93 88.04 90.22 88.33 ;
      RECT  90.38 85.44 90.7 85.76 ;
      RECT  89.19 85.92 89.52 86.07 ;
      RECT  89.87 85.44 90.19 85.76 ;
      RECT  90.35 88.58 90.64 88.87 ;
      RECT  89.01 89.94 91.61 90.23 ;
      RECT  89.21 86.07 89.5 86.23 ;
      RECT  89.01 84.86 91.61 85.15 ;
      RECT  89.93 92.14 90.22 91.85 ;
      RECT  90.38 94.74 90.7 94.42 ;
      RECT  89.19 94.26 89.52 94.11 ;
      RECT  89.87 94.74 90.19 94.42 ;
      RECT  90.35 91.6 90.64 91.31 ;
      RECT  89.01 90.24 91.61 89.95 ;
      RECT  89.21 94.11 89.5 93.95 ;
      RECT  89.01 95.32 91.61 95.03 ;
      RECT  89.93 98.22 90.22 98.51 ;
      RECT  90.38 95.62 90.7 95.94 ;
      RECT  89.19 96.1 89.52 96.25 ;
      RECT  89.87 95.62 90.19 95.94 ;
      RECT  90.35 98.76 90.64 99.05 ;
      RECT  89.01 100.12 91.61 100.41 ;
      RECT  89.21 96.25 89.5 96.41 ;
      RECT  89.01 95.04 91.61 95.33 ;
      RECT  89.93 102.32 90.22 102.03 ;
      RECT  90.38 104.92 90.7 104.6 ;
      RECT  89.19 104.44 89.52 104.29 ;
      RECT  89.87 104.92 90.19 104.6 ;
      RECT  90.35 101.78 90.64 101.49 ;
      RECT  89.01 100.42 91.61 100.13 ;
      RECT  89.21 104.29 89.5 104.13 ;
      RECT  89.01 105.5 91.61 105.21 ;
      RECT  89.93 108.4 90.22 108.69 ;
      RECT  90.38 105.8 90.7 106.12 ;
      RECT  89.19 106.28 89.52 106.43 ;
      RECT  89.87 105.8 90.19 106.12 ;
      RECT  90.35 108.94 90.64 109.23 ;
      RECT  89.01 110.3 91.61 110.59 ;
      RECT  89.21 106.43 89.5 106.59 ;
      RECT  89.01 105.22 91.61 105.51 ;
      RECT  89.93 112.5 90.22 112.21 ;
      RECT  90.38 115.1 90.7 114.78 ;
      RECT  89.19 114.62 89.52 114.47 ;
      RECT  89.87 115.1 90.19 114.78 ;
      RECT  90.35 111.96 90.64 111.67 ;
      RECT  89.01 110.6 91.61 110.31 ;
      RECT  89.21 114.47 89.5 114.31 ;
      RECT  89.01 115.68 91.61 115.39 ;
      RECT  89.93 118.58 90.22 118.87 ;
      RECT  90.38 115.98 90.7 116.3 ;
      RECT  89.19 116.46 89.52 116.61 ;
      RECT  89.87 115.98 90.19 116.3 ;
      RECT  90.35 119.12 90.64 119.41 ;
      RECT  89.01 120.48 91.61 120.77 ;
      RECT  89.21 116.61 89.5 116.77 ;
      RECT  89.01 115.4 91.61 115.69 ;
      RECT  89.01 24.99 91.61 25.15 ;
      RECT  89.01 32.87 91.61 33.03 ;
      RECT  89.01 35.17 91.61 35.33 ;
      RECT  89.01 43.05 91.61 43.21 ;
      RECT  89.01 45.35 91.61 45.51 ;
      RECT  89.01 53.23 91.61 53.39 ;
      RECT  89.01 55.53 91.61 55.69 ;
      RECT  89.01 63.41 91.61 63.57 ;
      RECT  89.01 65.71 91.61 65.87 ;
      RECT  89.01 73.59 91.61 73.75 ;
      RECT  89.01 75.89 91.61 76.05 ;
      RECT  89.01 83.77 91.61 83.93 ;
      RECT  89.01 86.07 91.61 86.23 ;
      RECT  89.01 93.95 91.61 94.11 ;
      RECT  89.01 96.25 91.61 96.41 ;
      RECT  89.01 104.13 91.61 104.29 ;
      RECT  89.01 106.43 91.61 106.59 ;
      RECT  89.01 114.31 91.61 114.47 ;
      RECT  89.01 116.61 91.61 116.77 ;
      RECT  89.01 100.13 91.61 100.42 ;
      RECT  89.01 79.77 91.61 80.06 ;
      RECT  89.01 69.58 91.61 69.87 ;
      RECT  89.01 69.59 91.61 69.88 ;
      RECT  89.01 49.22 91.61 49.51 ;
      RECT  89.01 100.12 91.61 100.41 ;
      RECT  89.01 39.05 91.61 39.34 ;
      RECT  89.01 89.94 91.61 90.23 ;
      RECT  89.01 110.31 91.61 110.6 ;
      RECT  89.01 89.95 91.61 90.24 ;
      RECT  89.01 39.04 91.61 39.33 ;
      RECT  89.01 59.4 91.61 59.69 ;
      RECT  89.01 59.41 91.61 59.7 ;
      RECT  89.01 110.3 91.61 110.59 ;
      RECT  89.01 28.87 91.61 29.16 ;
      RECT  89.01 49.23 91.61 49.52 ;
      RECT  89.01 79.76 91.61 80.05 ;
      RECT  89.01 64.5 91.61 64.79 ;
      RECT  89.01 115.39 91.61 115.68 ;
      RECT  89.01 64.49 91.61 64.78 ;
      RECT  89.01 95.03 91.61 95.32 ;
      RECT  89.01 33.96 91.61 34.25 ;
      RECT  89.01 44.14 91.61 44.43 ;
      RECT  89.01 84.85 91.61 85.14 ;
      RECT  89.01 54.31 91.61 54.6 ;
      RECT  89.01 105.22 91.61 105.51 ;
      RECT  89.01 105.21 91.61 105.5 ;
      RECT  89.01 54.32 91.61 54.61 ;
      RECT  89.01 44.13 91.61 44.42 ;
      RECT  89.01 95.04 91.61 95.33 ;
      RECT  89.01 74.67 91.61 74.96 ;
      RECT  89.01 74.68 91.61 74.97 ;
      RECT  89.01 33.95 91.61 34.24 ;
      RECT  89.01 84.86 91.61 85.15 ;
      RECT  92.53 31.06 92.82 30.77 ;
      RECT  92.98 33.66 93.3 33.34 ;
      RECT  91.79 33.18 92.12 33.03 ;
      RECT  92.47 33.66 92.79 33.34 ;
      RECT  92.95 30.52 93.24 30.23 ;
      RECT  91.61 29.16 94.21 28.87 ;
      RECT  91.81 33.03 92.1 32.87 ;
      RECT  91.61 34.24 94.21 33.95 ;
      RECT  95.13 31.06 95.42 30.77 ;
      RECT  95.58 33.66 95.9 33.34 ;
      RECT  94.39 33.18 94.72 33.03 ;
      RECT  95.07 33.66 95.39 33.34 ;
      RECT  95.55 30.52 95.84 30.23 ;
      RECT  94.21 29.16 96.81 28.87 ;
      RECT  94.41 33.03 94.7 32.87 ;
      RECT  94.21 34.24 96.81 33.95 ;
      RECT  91.61 33.03 96.81 32.87 ;
      RECT  94.21 29.16 96.81 28.87 ;
      RECT  91.61 29.16 94.21 28.87 ;
      RECT  91.61 34.24 94.21 33.95 ;
      RECT  94.21 34.24 96.81 33.95 ;
      RECT  92.53 26.96 92.82 27.25 ;
      RECT  92.98 24.36 93.3 24.68 ;
      RECT  91.79 24.84 92.12 24.99 ;
      RECT  92.47 24.36 92.79 24.68 ;
      RECT  92.95 27.5 93.24 27.79 ;
      RECT  91.61 28.86 94.21 29.15 ;
      RECT  91.81 24.99 92.1 25.15 ;
      RECT  91.61 23.78 94.21 24.07 ;
      RECT  95.13 26.96 95.42 27.25 ;
      RECT  95.58 24.36 95.9 24.68 ;
      RECT  94.39 24.84 94.72 24.99 ;
      RECT  95.07 24.36 95.39 24.68 ;
      RECT  95.55 27.5 95.84 27.79 ;
      RECT  94.21 28.86 96.81 29.15 ;
      RECT  94.41 24.99 94.7 25.15 ;
      RECT  94.21 23.78 96.81 24.07 ;
      RECT  91.61 24.99 96.81 25.15 ;
      RECT  94.21 28.86 96.81 29.15 ;
      RECT  91.61 28.86 94.21 29.15 ;
      RECT  91.61 23.78 94.21 24.07 ;
      RECT  94.21 23.78 96.81 24.07 ;
      RECT  92.53 118.58 92.82 118.87 ;
      RECT  92.98 115.98 93.3 116.3 ;
      RECT  91.79 116.46 92.12 116.61 ;
      RECT  92.47 115.98 92.79 116.3 ;
      RECT  92.95 119.12 93.24 119.41 ;
      RECT  91.61 120.48 94.21 120.77 ;
      RECT  91.81 116.61 92.1 116.77 ;
      RECT  91.61 115.4 94.21 115.69 ;
      RECT  95.13 118.58 95.42 118.87 ;
      RECT  95.58 115.98 95.9 116.3 ;
      RECT  94.39 116.46 94.72 116.61 ;
      RECT  95.07 115.98 95.39 116.3 ;
      RECT  95.55 119.12 95.84 119.41 ;
      RECT  94.21 120.48 96.81 120.77 ;
      RECT  94.41 116.61 94.7 116.77 ;
      RECT  94.21 115.4 96.81 115.69 ;
      RECT  91.61 116.61 96.81 116.77 ;
      RECT  94.21 120.48 96.81 120.77 ;
      RECT  91.61 120.48 94.21 120.77 ;
      RECT  91.61 115.4 94.21 115.69 ;
      RECT  94.21 115.4 96.81 115.69 ;
      RECT  87.33 26.96 87.62 27.25 ;
      RECT  87.78 24.36 88.1 24.68 ;
      RECT  86.59 24.84 86.92 24.99 ;
      RECT  87.27 24.36 87.59 24.68 ;
      RECT  87.75 27.5 88.04 27.79 ;
      RECT  86.41 28.86 89.01 29.15 ;
      RECT  86.61 24.99 86.9 25.15 ;
      RECT  86.41 23.78 89.01 24.07 ;
      RECT  87.33 31.06 87.62 30.77 ;
      RECT  87.78 33.66 88.1 33.34 ;
      RECT  86.59 33.18 86.92 33.03 ;
      RECT  87.27 33.66 87.59 33.34 ;
      RECT  87.75 30.52 88.04 30.23 ;
      RECT  86.41 29.16 89.01 28.87 ;
      RECT  86.61 33.03 86.9 32.87 ;
      RECT  86.41 34.24 89.01 33.95 ;
      RECT  87.33 37.14 87.62 37.43 ;
      RECT  87.78 34.54 88.1 34.86 ;
      RECT  86.59 35.02 86.92 35.17 ;
      RECT  87.27 34.54 87.59 34.86 ;
      RECT  87.75 37.68 88.04 37.97 ;
      RECT  86.41 39.04 89.01 39.33 ;
      RECT  86.61 35.17 86.9 35.33 ;
      RECT  86.41 33.96 89.01 34.25 ;
      RECT  87.33 41.24 87.62 40.95 ;
      RECT  87.78 43.84 88.1 43.52 ;
      RECT  86.59 43.36 86.92 43.21 ;
      RECT  87.27 43.84 87.59 43.52 ;
      RECT  87.75 40.7 88.04 40.41 ;
      RECT  86.41 39.34 89.01 39.05 ;
      RECT  86.61 43.21 86.9 43.05 ;
      RECT  86.41 44.42 89.01 44.13 ;
      RECT  87.33 47.32 87.62 47.61 ;
      RECT  87.78 44.72 88.1 45.04 ;
      RECT  86.59 45.2 86.92 45.35 ;
      RECT  87.27 44.72 87.59 45.04 ;
      RECT  87.75 47.86 88.04 48.15 ;
      RECT  86.41 49.22 89.01 49.51 ;
      RECT  86.61 45.35 86.9 45.51 ;
      RECT  86.41 44.14 89.01 44.43 ;
      RECT  87.33 51.42 87.62 51.13 ;
      RECT  87.78 54.02 88.1 53.7 ;
      RECT  86.59 53.54 86.92 53.39 ;
      RECT  87.27 54.02 87.59 53.7 ;
      RECT  87.75 50.88 88.04 50.59 ;
      RECT  86.41 49.52 89.01 49.23 ;
      RECT  86.61 53.39 86.9 53.23 ;
      RECT  86.41 54.6 89.01 54.31 ;
      RECT  87.33 57.5 87.62 57.79 ;
      RECT  87.78 54.9 88.1 55.22 ;
      RECT  86.59 55.38 86.92 55.53 ;
      RECT  87.27 54.9 87.59 55.22 ;
      RECT  87.75 58.04 88.04 58.33 ;
      RECT  86.41 59.4 89.01 59.69 ;
      RECT  86.61 55.53 86.9 55.69 ;
      RECT  86.41 54.32 89.01 54.61 ;
      RECT  87.33 61.6 87.62 61.31 ;
      RECT  87.78 64.2 88.1 63.88 ;
      RECT  86.59 63.72 86.92 63.57 ;
      RECT  87.27 64.2 87.59 63.88 ;
      RECT  87.75 61.06 88.04 60.77 ;
      RECT  86.41 59.7 89.01 59.41 ;
      RECT  86.61 63.57 86.9 63.41 ;
      RECT  86.41 64.78 89.01 64.49 ;
      RECT  87.33 67.68 87.62 67.97 ;
      RECT  87.78 65.08 88.1 65.4 ;
      RECT  86.59 65.56 86.92 65.71 ;
      RECT  87.27 65.08 87.59 65.4 ;
      RECT  87.75 68.22 88.04 68.51 ;
      RECT  86.41 69.58 89.01 69.87 ;
      RECT  86.61 65.71 86.9 65.87 ;
      RECT  86.41 64.5 89.01 64.79 ;
      RECT  87.33 71.78 87.62 71.49 ;
      RECT  87.78 74.38 88.1 74.06 ;
      RECT  86.59 73.9 86.92 73.75 ;
      RECT  87.27 74.38 87.59 74.06 ;
      RECT  87.75 71.24 88.04 70.95 ;
      RECT  86.41 69.88 89.01 69.59 ;
      RECT  86.61 73.75 86.9 73.59 ;
      RECT  86.41 74.96 89.01 74.67 ;
      RECT  87.33 77.86 87.62 78.15 ;
      RECT  87.78 75.26 88.1 75.58 ;
      RECT  86.59 75.74 86.92 75.89 ;
      RECT  87.27 75.26 87.59 75.58 ;
      RECT  87.75 78.4 88.04 78.69 ;
      RECT  86.41 79.76 89.01 80.05 ;
      RECT  86.61 75.89 86.9 76.05 ;
      RECT  86.41 74.68 89.01 74.97 ;
      RECT  87.33 81.96 87.62 81.67 ;
      RECT  87.78 84.56 88.1 84.24 ;
      RECT  86.59 84.08 86.92 83.93 ;
      RECT  87.27 84.56 87.59 84.24 ;
      RECT  87.75 81.42 88.04 81.13 ;
      RECT  86.41 80.06 89.01 79.77 ;
      RECT  86.61 83.93 86.9 83.77 ;
      RECT  86.41 85.14 89.01 84.85 ;
      RECT  87.33 88.04 87.62 88.33 ;
      RECT  87.78 85.44 88.1 85.76 ;
      RECT  86.59 85.92 86.92 86.07 ;
      RECT  87.27 85.44 87.59 85.76 ;
      RECT  87.75 88.58 88.04 88.87 ;
      RECT  86.41 89.94 89.01 90.23 ;
      RECT  86.61 86.07 86.9 86.23 ;
      RECT  86.41 84.86 89.01 85.15 ;
      RECT  87.33 92.14 87.62 91.85 ;
      RECT  87.78 94.74 88.1 94.42 ;
      RECT  86.59 94.26 86.92 94.11 ;
      RECT  87.27 94.74 87.59 94.42 ;
      RECT  87.75 91.6 88.04 91.31 ;
      RECT  86.41 90.24 89.01 89.95 ;
      RECT  86.61 94.11 86.9 93.95 ;
      RECT  86.41 95.32 89.01 95.03 ;
      RECT  87.33 98.22 87.62 98.51 ;
      RECT  87.78 95.62 88.1 95.94 ;
      RECT  86.59 96.1 86.92 96.25 ;
      RECT  87.27 95.62 87.59 95.94 ;
      RECT  87.75 98.76 88.04 99.05 ;
      RECT  86.41 100.12 89.01 100.41 ;
      RECT  86.61 96.25 86.9 96.41 ;
      RECT  86.41 95.04 89.01 95.33 ;
      RECT  87.33 102.32 87.62 102.03 ;
      RECT  87.78 104.92 88.1 104.6 ;
      RECT  86.59 104.44 86.92 104.29 ;
      RECT  87.27 104.92 87.59 104.6 ;
      RECT  87.75 101.78 88.04 101.49 ;
      RECT  86.41 100.42 89.01 100.13 ;
      RECT  86.61 104.29 86.9 104.13 ;
      RECT  86.41 105.5 89.01 105.21 ;
      RECT  87.33 108.4 87.62 108.69 ;
      RECT  87.78 105.8 88.1 106.12 ;
      RECT  86.59 106.28 86.92 106.43 ;
      RECT  87.27 105.8 87.59 106.12 ;
      RECT  87.75 108.94 88.04 109.23 ;
      RECT  86.41 110.3 89.01 110.59 ;
      RECT  86.61 106.43 86.9 106.59 ;
      RECT  86.41 105.22 89.01 105.51 ;
      RECT  87.33 112.5 87.62 112.21 ;
      RECT  87.78 115.1 88.1 114.78 ;
      RECT  86.59 114.62 86.92 114.47 ;
      RECT  87.27 115.1 87.59 114.78 ;
      RECT  87.75 111.96 88.04 111.67 ;
      RECT  86.41 110.6 89.01 110.31 ;
      RECT  86.61 114.47 86.9 114.31 ;
      RECT  86.41 115.68 89.01 115.39 ;
      RECT  87.33 118.58 87.62 118.87 ;
      RECT  87.78 115.98 88.1 116.3 ;
      RECT  86.59 116.46 86.92 116.61 ;
      RECT  87.27 115.98 87.59 116.3 ;
      RECT  87.75 119.12 88.04 119.41 ;
      RECT  86.41 120.48 89.01 120.77 ;
      RECT  86.61 116.61 86.9 116.77 ;
      RECT  86.41 115.4 89.01 115.69 ;
      RECT  86.41 24.99 89.01 25.15 ;
      RECT  86.41 32.87 89.01 33.03 ;
      RECT  86.41 35.17 89.01 35.33 ;
      RECT  86.41 43.05 89.01 43.21 ;
      RECT  86.41 45.35 89.01 45.51 ;
      RECT  86.41 53.23 89.01 53.39 ;
      RECT  86.41 55.53 89.01 55.69 ;
      RECT  86.41 63.41 89.01 63.57 ;
      RECT  86.41 65.71 89.01 65.87 ;
      RECT  86.41 73.59 89.01 73.75 ;
      RECT  86.41 75.89 89.01 76.05 ;
      RECT  86.41 83.77 89.01 83.93 ;
      RECT  86.41 86.07 89.01 86.23 ;
      RECT  86.41 93.95 89.01 94.11 ;
      RECT  86.41 96.25 89.01 96.41 ;
      RECT  86.41 104.13 89.01 104.29 ;
      RECT  86.41 106.43 89.01 106.59 ;
      RECT  86.41 114.31 89.01 114.47 ;
      RECT  86.41 116.61 89.01 116.77 ;
      RECT  86.41 100.13 89.01 100.42 ;
      RECT  86.41 79.77 89.01 80.06 ;
      RECT  86.41 69.58 89.01 69.87 ;
      RECT  86.41 69.59 89.01 69.88 ;
      RECT  86.41 49.22 89.01 49.51 ;
      RECT  86.41 100.12 89.01 100.41 ;
      RECT  86.41 39.05 89.01 39.34 ;
      RECT  86.41 89.94 89.01 90.23 ;
      RECT  86.41 120.48 89.01 120.77 ;
      RECT  86.41 110.31 89.01 110.6 ;
      RECT  86.41 89.95 89.01 90.24 ;
      RECT  86.41 39.04 89.01 39.33 ;
      RECT  86.41 59.4 89.01 59.69 ;
      RECT  86.41 59.41 89.01 59.7 ;
      RECT  86.41 28.86 89.01 29.15 ;
      RECT  86.41 110.3 89.01 110.59 ;
      RECT  86.41 28.87 89.01 29.16 ;
      RECT  86.41 49.23 89.01 49.52 ;
      RECT  86.41 79.76 89.01 80.05 ;
      RECT  86.41 64.5 89.01 64.79 ;
      RECT  86.41 115.39 89.01 115.68 ;
      RECT  86.41 64.49 89.01 64.78 ;
      RECT  86.41 95.03 89.01 95.32 ;
      RECT  86.41 23.78 89.01 24.07 ;
      RECT  86.41 115.4 89.01 115.69 ;
      RECT  86.41 33.96 89.01 34.25 ;
      RECT  86.41 44.14 89.01 44.43 ;
      RECT  86.41 84.85 89.01 85.14 ;
      RECT  86.41 54.31 89.01 54.6 ;
      RECT  86.41 105.22 89.01 105.51 ;
      RECT  86.41 105.21 89.01 105.5 ;
      RECT  86.41 54.32 89.01 54.61 ;
      RECT  86.41 44.13 89.01 44.42 ;
      RECT  86.41 95.04 89.01 95.33 ;
      RECT  86.41 74.67 89.01 74.96 ;
      RECT  86.41 74.68 89.01 74.97 ;
      RECT  86.41 33.95 89.01 34.24 ;
      RECT  86.41 84.86 89.01 85.15 ;
      RECT  97.73 26.96 98.02 27.25 ;
      RECT  98.18 24.36 98.5 24.68 ;
      RECT  96.99 24.84 97.32 24.99 ;
      RECT  97.67 24.36 97.99 24.68 ;
      RECT  98.15 27.5 98.44 27.79 ;
      RECT  96.81 28.86 99.41 29.15 ;
      RECT  97.01 24.99 97.3 25.15 ;
      RECT  96.81 23.78 99.41 24.07 ;
      RECT  97.73 31.06 98.02 30.77 ;
      RECT  98.18 33.66 98.5 33.34 ;
      RECT  96.99 33.18 97.32 33.03 ;
      RECT  97.67 33.66 97.99 33.34 ;
      RECT  98.15 30.52 98.44 30.23 ;
      RECT  96.81 29.16 99.41 28.87 ;
      RECT  97.01 33.03 97.3 32.87 ;
      RECT  96.81 34.24 99.41 33.95 ;
      RECT  97.73 37.14 98.02 37.43 ;
      RECT  98.18 34.54 98.5 34.86 ;
      RECT  96.99 35.02 97.32 35.17 ;
      RECT  97.67 34.54 97.99 34.86 ;
      RECT  98.15 37.68 98.44 37.97 ;
      RECT  96.81 39.04 99.41 39.33 ;
      RECT  97.01 35.17 97.3 35.33 ;
      RECT  96.81 33.96 99.41 34.25 ;
      RECT  97.73 41.24 98.02 40.95 ;
      RECT  98.18 43.84 98.5 43.52 ;
      RECT  96.99 43.36 97.32 43.21 ;
      RECT  97.67 43.84 97.99 43.52 ;
      RECT  98.15 40.7 98.44 40.41 ;
      RECT  96.81 39.34 99.41 39.05 ;
      RECT  97.01 43.21 97.3 43.05 ;
      RECT  96.81 44.42 99.41 44.13 ;
      RECT  97.73 47.32 98.02 47.61 ;
      RECT  98.18 44.72 98.5 45.04 ;
      RECT  96.99 45.2 97.32 45.35 ;
      RECT  97.67 44.72 97.99 45.04 ;
      RECT  98.15 47.86 98.44 48.15 ;
      RECT  96.81 49.22 99.41 49.51 ;
      RECT  97.01 45.35 97.3 45.51 ;
      RECT  96.81 44.14 99.41 44.43 ;
      RECT  97.73 51.42 98.02 51.13 ;
      RECT  98.18 54.02 98.5 53.7 ;
      RECT  96.99 53.54 97.32 53.39 ;
      RECT  97.67 54.02 97.99 53.7 ;
      RECT  98.15 50.88 98.44 50.59 ;
      RECT  96.81 49.52 99.41 49.23 ;
      RECT  97.01 53.39 97.3 53.23 ;
      RECT  96.81 54.6 99.41 54.31 ;
      RECT  97.73 57.5 98.02 57.79 ;
      RECT  98.18 54.9 98.5 55.22 ;
      RECT  96.99 55.38 97.32 55.53 ;
      RECT  97.67 54.9 97.99 55.22 ;
      RECT  98.15 58.04 98.44 58.33 ;
      RECT  96.81 59.4 99.41 59.69 ;
      RECT  97.01 55.53 97.3 55.69 ;
      RECT  96.81 54.32 99.41 54.61 ;
      RECT  97.73 61.6 98.02 61.31 ;
      RECT  98.18 64.2 98.5 63.88 ;
      RECT  96.99 63.72 97.32 63.57 ;
      RECT  97.67 64.2 97.99 63.88 ;
      RECT  98.15 61.06 98.44 60.77 ;
      RECT  96.81 59.7 99.41 59.41 ;
      RECT  97.01 63.57 97.3 63.41 ;
      RECT  96.81 64.78 99.41 64.49 ;
      RECT  97.73 67.68 98.02 67.97 ;
      RECT  98.18 65.08 98.5 65.4 ;
      RECT  96.99 65.56 97.32 65.71 ;
      RECT  97.67 65.08 97.99 65.4 ;
      RECT  98.15 68.22 98.44 68.51 ;
      RECT  96.81 69.58 99.41 69.87 ;
      RECT  97.01 65.71 97.3 65.87 ;
      RECT  96.81 64.5 99.41 64.79 ;
      RECT  97.73 71.78 98.02 71.49 ;
      RECT  98.18 74.38 98.5 74.06 ;
      RECT  96.99 73.9 97.32 73.75 ;
      RECT  97.67 74.38 97.99 74.06 ;
      RECT  98.15 71.24 98.44 70.95 ;
      RECT  96.81 69.88 99.41 69.59 ;
      RECT  97.01 73.75 97.3 73.59 ;
      RECT  96.81 74.96 99.41 74.67 ;
      RECT  97.73 77.86 98.02 78.15 ;
      RECT  98.18 75.26 98.5 75.58 ;
      RECT  96.99 75.74 97.32 75.89 ;
      RECT  97.67 75.26 97.99 75.58 ;
      RECT  98.15 78.4 98.44 78.69 ;
      RECT  96.81 79.76 99.41 80.05 ;
      RECT  97.01 75.89 97.3 76.05 ;
      RECT  96.81 74.68 99.41 74.97 ;
      RECT  97.73 81.96 98.02 81.67 ;
      RECT  98.18 84.56 98.5 84.24 ;
      RECT  96.99 84.08 97.32 83.93 ;
      RECT  97.67 84.56 97.99 84.24 ;
      RECT  98.15 81.42 98.44 81.13 ;
      RECT  96.81 80.06 99.41 79.77 ;
      RECT  97.01 83.93 97.3 83.77 ;
      RECT  96.81 85.14 99.41 84.85 ;
      RECT  97.73 88.04 98.02 88.33 ;
      RECT  98.18 85.44 98.5 85.76 ;
      RECT  96.99 85.92 97.32 86.07 ;
      RECT  97.67 85.44 97.99 85.76 ;
      RECT  98.15 88.58 98.44 88.87 ;
      RECT  96.81 89.94 99.41 90.23 ;
      RECT  97.01 86.07 97.3 86.23 ;
      RECT  96.81 84.86 99.41 85.15 ;
      RECT  97.73 92.14 98.02 91.85 ;
      RECT  98.18 94.74 98.5 94.42 ;
      RECT  96.99 94.26 97.32 94.11 ;
      RECT  97.67 94.74 97.99 94.42 ;
      RECT  98.15 91.6 98.44 91.31 ;
      RECT  96.81 90.24 99.41 89.95 ;
      RECT  97.01 94.11 97.3 93.95 ;
      RECT  96.81 95.32 99.41 95.03 ;
      RECT  97.73 98.22 98.02 98.51 ;
      RECT  98.18 95.62 98.5 95.94 ;
      RECT  96.99 96.1 97.32 96.25 ;
      RECT  97.67 95.62 97.99 95.94 ;
      RECT  98.15 98.76 98.44 99.05 ;
      RECT  96.81 100.12 99.41 100.41 ;
      RECT  97.01 96.25 97.3 96.41 ;
      RECT  96.81 95.04 99.41 95.33 ;
      RECT  97.73 102.32 98.02 102.03 ;
      RECT  98.18 104.92 98.5 104.6 ;
      RECT  96.99 104.44 97.32 104.29 ;
      RECT  97.67 104.92 97.99 104.6 ;
      RECT  98.15 101.78 98.44 101.49 ;
      RECT  96.81 100.42 99.41 100.13 ;
      RECT  97.01 104.29 97.3 104.13 ;
      RECT  96.81 105.5 99.41 105.21 ;
      RECT  97.73 108.4 98.02 108.69 ;
      RECT  98.18 105.8 98.5 106.12 ;
      RECT  96.99 106.28 97.32 106.43 ;
      RECT  97.67 105.8 97.99 106.12 ;
      RECT  98.15 108.94 98.44 109.23 ;
      RECT  96.81 110.3 99.41 110.59 ;
      RECT  97.01 106.43 97.3 106.59 ;
      RECT  96.81 105.22 99.41 105.51 ;
      RECT  97.73 112.5 98.02 112.21 ;
      RECT  98.18 115.1 98.5 114.78 ;
      RECT  96.99 114.62 97.32 114.47 ;
      RECT  97.67 115.1 97.99 114.78 ;
      RECT  98.15 111.96 98.44 111.67 ;
      RECT  96.81 110.6 99.41 110.31 ;
      RECT  97.01 114.47 97.3 114.31 ;
      RECT  96.81 115.68 99.41 115.39 ;
      RECT  97.73 118.58 98.02 118.87 ;
      RECT  98.18 115.98 98.5 116.3 ;
      RECT  96.99 116.46 97.32 116.61 ;
      RECT  97.67 115.98 97.99 116.3 ;
      RECT  98.15 119.12 98.44 119.41 ;
      RECT  96.81 120.48 99.41 120.77 ;
      RECT  97.01 116.61 97.3 116.77 ;
      RECT  96.81 115.4 99.41 115.69 ;
      RECT  96.81 24.99 99.41 25.15 ;
      RECT  96.81 32.87 99.41 33.03 ;
      RECT  96.81 35.17 99.41 35.33 ;
      RECT  96.81 43.05 99.41 43.21 ;
      RECT  96.81 45.35 99.41 45.51 ;
      RECT  96.81 53.23 99.41 53.39 ;
      RECT  96.81 55.53 99.41 55.69 ;
      RECT  96.81 63.41 99.41 63.57 ;
      RECT  96.81 65.71 99.41 65.87 ;
      RECT  96.81 73.59 99.41 73.75 ;
      RECT  96.81 75.89 99.41 76.05 ;
      RECT  96.81 83.77 99.41 83.93 ;
      RECT  96.81 86.07 99.41 86.23 ;
      RECT  96.81 93.95 99.41 94.11 ;
      RECT  96.81 96.25 99.41 96.41 ;
      RECT  96.81 104.13 99.41 104.29 ;
      RECT  96.81 106.43 99.41 106.59 ;
      RECT  96.81 114.31 99.41 114.47 ;
      RECT  96.81 116.61 99.41 116.77 ;
      RECT  96.81 100.13 99.41 100.42 ;
      RECT  96.81 79.77 99.41 80.06 ;
      RECT  96.81 69.58 99.41 69.87 ;
      RECT  96.81 69.59 99.41 69.88 ;
      RECT  96.81 49.22 99.41 49.51 ;
      RECT  96.81 100.12 99.41 100.41 ;
      RECT  96.81 39.05 99.41 39.34 ;
      RECT  96.81 89.94 99.41 90.23 ;
      RECT  96.81 120.48 99.41 120.77 ;
      RECT  96.81 110.31 99.41 110.6 ;
      RECT  96.81 89.95 99.41 90.24 ;
      RECT  96.81 39.04 99.41 39.33 ;
      RECT  96.81 59.4 99.41 59.69 ;
      RECT  96.81 59.41 99.41 59.7 ;
      RECT  96.81 28.86 99.41 29.15 ;
      RECT  96.81 110.3 99.41 110.59 ;
      RECT  96.81 28.87 99.41 29.16 ;
      RECT  96.81 49.23 99.41 49.52 ;
      RECT  96.81 79.76 99.41 80.05 ;
      RECT  96.81 64.5 99.41 64.79 ;
      RECT  96.81 115.39 99.41 115.68 ;
      RECT  96.81 64.49 99.41 64.78 ;
      RECT  96.81 95.03 99.41 95.32 ;
      RECT  96.81 23.78 99.41 24.07 ;
      RECT  96.81 115.4 99.41 115.69 ;
      RECT  96.81 33.96 99.41 34.25 ;
      RECT  96.81 44.14 99.41 44.43 ;
      RECT  96.81 84.85 99.41 85.14 ;
      RECT  96.81 54.31 99.41 54.6 ;
      RECT  96.81 105.22 99.41 105.51 ;
      RECT  96.81 105.21 99.41 105.5 ;
      RECT  96.81 54.32 99.41 54.61 ;
      RECT  96.81 44.13 99.41 44.42 ;
      RECT  96.81 95.04 99.41 95.33 ;
      RECT  96.81 74.67 99.41 74.96 ;
      RECT  96.81 74.68 99.41 74.97 ;
      RECT  96.81 33.95 99.41 34.24 ;
      RECT  96.81 84.86 99.41 85.15 ;
      RECT  85.72 32.87 100.1 33.03 ;
      RECT  85.72 35.17 100.1 35.33 ;
      RECT  85.72 43.05 100.1 43.21 ;
      RECT  85.72 45.35 100.1 45.51 ;
      RECT  85.72 53.23 100.1 53.39 ;
      RECT  85.72 55.53 100.1 55.69 ;
      RECT  85.72 63.41 100.1 63.57 ;
      RECT  85.72 65.71 100.1 65.87 ;
      RECT  85.72 73.59 100.1 73.75 ;
      RECT  85.72 75.89 100.1 76.05 ;
      RECT  85.72 83.77 100.1 83.93 ;
      RECT  85.72 86.07 100.1 86.23 ;
      RECT  85.72 93.95 100.1 94.11 ;
      RECT  85.72 96.25 100.1 96.41 ;
      RECT  85.72 104.13 100.1 104.29 ;
      RECT  85.72 106.43 100.1 106.59 ;
      RECT  85.72 114.31 100.1 114.47 ;
      RECT  89.01 39.04 91.61 39.33 ;
      RECT  89.01 69.59 91.61 69.88 ;
      RECT  89.01 59.41 91.61 59.7 ;
      RECT  89.01 89.94 91.61 90.23 ;
      RECT  89.01 69.58 91.61 69.87 ;
      RECT  89.01 49.23 91.61 49.52 ;
      RECT  89.01 28.87 91.61 29.16 ;
      RECT  89.01 59.4 91.61 59.69 ;
      RECT  89.01 49.22 91.61 49.51 ;
      RECT  89.01 100.12 91.61 100.41 ;
      RECT  89.01 110.3 91.61 110.59 ;
      RECT  89.01 79.77 91.61 80.06 ;
      RECT  89.01 100.13 91.61 100.42 ;
      RECT  89.01 79.76 91.61 80.05 ;
      RECT  89.01 39.05 91.61 39.34 ;
      RECT  89.01 110.31 91.61 110.6 ;
      RECT  89.01 89.95 91.61 90.24 ;
      RECT  89.01 54.31 91.61 54.6 ;
      RECT  89.01 64.49 91.61 64.78 ;
      RECT  89.01 84.85 91.61 85.14 ;
      RECT  89.01 44.13 91.61 44.42 ;
      RECT  89.01 105.22 91.61 105.51 ;
      RECT  89.01 44.14 91.61 44.43 ;
      RECT  89.01 84.86 91.61 85.15 ;
      RECT  89.01 115.39 91.61 115.68 ;
      RECT  89.01 74.67 91.61 74.96 ;
      RECT  89.01 64.5 91.61 64.79 ;
      RECT  89.01 95.04 91.61 95.33 ;
      RECT  89.01 74.68 91.61 74.97 ;
      RECT  89.01 54.32 91.61 54.61 ;
      RECT  89.01 95.03 91.61 95.32 ;
      RECT  89.01 105.21 91.61 105.5 ;
      RECT  89.01 33.96 91.61 34.25 ;
      RECT  89.01 33.95 91.61 34.24 ;
      RECT  89.01 14.37 91.61 14.51 ;
      RECT  91.61 14.37 94.21 14.51 ;
      RECT  94.21 14.37 96.81 14.51 ;
      RECT  85.72 14.37 96.81 14.51 ;
      RECT  91.78 10.15 95.05 10.44 ;
      RECT  92.96 9.19 93.29 9.83 ;
      RECT  96.05 9.45 97.38 9.78 ;
      RECT  91.31 12.59 97.38 12.92 ;
      RECT  91.31 9.17 91.65 9.83 ;
      RECT  91.31 8.22 97.38 8.55 ;
      RECT  96.9 10.12 97.23 10.72 ;
      RECT  94.38 10.15 97.65 10.44 ;
      RECT  95.56 9.19 95.89 9.83 ;
      RECT  98.65 9.45 99.98 9.78 ;
      RECT  93.91 12.59 99.98 12.92 ;
      RECT  93.91 9.17 94.25 9.83 ;
      RECT  93.91 8.22 99.98 8.55 ;
      RECT  99.5 10.12 99.83 10.72 ;
      RECT  85.72 9.54 99.98 9.68 ;
      RECT  94.38 3.55 94.68 3.6 ;
      RECT  92.78 6.94 105.02 7.39 ;
      RECT  92.78 1.19 105.02 1.52 ;
      RECT  94.38 3.8 94.68 3.85 ;
      RECT  102.55 3.97 102.88 4.01 ;
      RECT  96.69 3.08 96.99 5.7 ;
      RECT  103.0 5.41 103.3 5.7 ;
      RECT  103.04 3.37 103.3 5.41 ;
      RECT  103.0 3.08 103.3 3.37 ;
      RECT  104.55 4.41 104.85 4.7 ;
      RECT  104.71 3.04 105.01 3.33 ;
      RECT  92.78 3.6 94.68 3.8 ;
      RECT  92.88 3.02 93.21 3.35 ;
      RECT  97.94 3.68 102.88 3.97 ;
      RECT  98.39 4.41 102.22 4.7 ;
      RECT  96.98 3.55 97.28 3.6 ;
      RECT  95.38 6.94 107.62 7.39 ;
      RECT  95.38 1.19 107.62 1.52 ;
      RECT  96.98 3.8 97.28 3.85 ;
      RECT  105.15 3.97 105.48 4.01 ;
      RECT  99.29 3.08 99.59 5.7 ;
      RECT  105.6 5.41 105.9 5.7 ;
      RECT  105.64 3.37 105.9 5.41 ;
      RECT  105.6 3.08 105.9 3.37 ;
      RECT  107.15 4.41 107.45 4.7 ;
      RECT  107.31 3.04 107.61 3.33 ;
      RECT  95.38 3.6 97.28 3.8 ;
      RECT  95.48 3.02 95.81 3.35 ;
      RECT  100.54 3.68 105.48 3.97 ;
      RECT  100.99 4.41 104.82 4.7 ;
      RECT  85.72 3.68 107.62 3.82 ;
      RECT  85.72 9.68 99.98 9.54 ;
      RECT  85.72 14.51 96.81 14.37 ;
      RECT  85.72 3.82 107.62 3.68 ;
      RECT  -100.18 -7.14 -99.85 -7.13 ;
      RECT  -102.42 -8.08 -100.97 -7.88 ;
      RECT  -100.18 -7.38 -99.85 -7.35 ;
      RECT  -94.38 -7.14 -94.05 -7.13 ;
      RECT  -102.42 -7.88 -102.13 -7.82 ;
      RECT  -93.24 -7.48 -92.61 -7.16 ;
      RECT  -95.46 -7.8 -95.26 -7.63 ;
      RECT  -95.46 -7.38 -95.26 -7.13 ;
      RECT  -94.77 -8.23 -91.24 -8.03 ;
      RECT  -100.18 -7.63 -95.26 -7.38 ;
      RECT  -101.26 -7.13 -95.77 -6.93 ;
      RECT  -101.3 -8.13 -100.97 -8.08 ;
      RECT  -103.29 -7.99 -102.61 -7.67 ;
      RECT  -96.1 -7.14 -95.77 -7.13 ;
      RECT  -101.3 -7.88 -100.97 -7.8 ;
      RECT  -103.31 -5.58 -90.66 -5.25 ;
      RECT  -91.58 -8.33 -91.24 -8.23 ;
      RECT  -100.18 -6.93 -99.85 -6.81 ;
      RECT  -91.58 -8.03 -91.24 -8.0 ;
      RECT  -101.26 -7.8 -101.06 -7.13 ;
      RECT  -95.46 -7.13 -94.05 -6.93 ;
      RECT  -96.1 -6.93 -95.77 -6.81 ;
      RECT  -95.5 -8.13 -95.17 -7.8 ;
      RECT  -100.57 -8.03 -100.27 -7.93 ;
      RECT  -97.61 -8.29 -97.28 -8.24 ;
      RECT  -103.37 -9.67 -90.84 -9.34 ;
      RECT  -102.14 -7.17 -101.51 -6.85 ;
      RECT  -100.57 -8.24 -97.28 -8.03 ;
      RECT  -94.77 -8.03 -94.47 -7.92 ;
      RECT  -94.38 -6.93 -94.05 -6.81 ;
      RECT  -100.18 -7.68 -99.85 -7.63 ;
      RECT  -97.61 -8.03 -97.28 -7.96 ;
      RECT  -102.42 -8.11 -102.13 -8.08 ;
      RECT  -103.31 -5.58 -66.43 -5.25 ;
      RECT  -103.37 -9.67 -66.49 -9.34 ;
      RECT  -100.18 -3.7 -99.85 -3.71 ;
      RECT  -102.42 -2.76 -100.97 -2.96 ;
      RECT  -100.18 -3.46 -99.85 -3.49 ;
      RECT  -94.38 -3.7 -94.05 -3.71 ;
      RECT  -102.42 -2.96 -102.13 -3.02 ;
      RECT  -93.24 -3.36 -92.61 -3.68 ;
      RECT  -95.46 -3.04 -95.26 -3.21 ;
      RECT  -95.46 -3.46 -95.26 -3.71 ;
      RECT  -94.77 -2.61 -91.24 -2.81 ;
      RECT  -100.18 -3.21 -95.26 -3.46 ;
      RECT  -101.26 -3.71 -95.77 -3.91 ;
      RECT  -101.3 -2.71 -100.97 -2.76 ;
      RECT  -103.29 -2.85 -102.61 -3.17 ;
      RECT  -96.1 -3.7 -95.77 -3.71 ;
      RECT  -101.3 -2.96 -100.97 -3.04 ;
      RECT  -103.31 -5.26 -90.66 -5.59 ;
      RECT  -91.58 -2.51 -91.24 -2.61 ;
      RECT  -100.18 -3.91 -99.85 -4.03 ;
      RECT  -91.58 -2.81 -91.24 -2.84 ;
      RECT  -101.26 -3.04 -101.06 -3.71 ;
      RECT  -95.46 -3.71 -94.05 -3.91 ;
      RECT  -96.1 -3.91 -95.77 -4.03 ;
      RECT  -95.5 -2.71 -95.17 -3.04 ;
      RECT  -100.57 -2.81 -100.27 -2.91 ;
      RECT  -97.61 -2.55 -97.28 -2.6 ;
      RECT  -103.37 -1.17 -90.84 -1.5 ;
      RECT  -102.14 -3.67 -101.51 -3.99 ;
      RECT  -100.57 -2.6 -97.28 -2.81 ;
      RECT  -94.77 -2.81 -94.47 -2.92 ;
      RECT  -94.38 -3.91 -94.05 -4.03 ;
      RECT  -100.18 -3.16 -99.85 -3.21 ;
      RECT  -97.61 -2.81 -97.28 -2.88 ;
      RECT  -102.42 -2.73 -102.13 -2.76 ;
      RECT  -103.31 -5.26 -66.43 -5.59 ;
      RECT  -103.37 -1.17 -66.49 -1.5 ;
      RECT  -10.54 85.14 -10.21 85.15 ;
      RECT  -12.78 84.2 -11.33 84.4 ;
      RECT  -10.54 84.9 -10.21 84.93 ;
      RECT  -4.74 85.14 -4.41 85.15 ;
      RECT  -12.78 84.4 -12.49 84.46 ;
      RECT  -3.6 84.8 -2.97 85.12 ;
      RECT  -5.82 84.48 -5.62 84.65 ;
      RECT  -5.82 84.9 -5.62 85.15 ;
      RECT  -5.13 84.05 -1.6 84.25 ;
      RECT  -10.54 84.65 -5.62 84.9 ;
      RECT  -11.62 85.15 -6.13 85.35 ;
      RECT  -11.66 84.15 -11.33 84.2 ;
      RECT  -13.65 84.29 -12.97 84.61 ;
      RECT  -6.46 85.14 -6.13 85.15 ;
      RECT  -11.66 84.4 -11.33 84.48 ;
      RECT  -13.67 86.7 -1.02 87.03 ;
      RECT  -1.94 83.95 -1.6 84.05 ;
      RECT  -10.54 85.35 -10.21 85.47 ;
      RECT  -1.94 84.25 -1.6 84.28 ;
      RECT  -11.62 84.48 -11.42 85.15 ;
      RECT  -5.82 85.15 -4.41 85.35 ;
      RECT  -6.46 85.35 -6.13 85.47 ;
      RECT  -5.86 84.15 -5.53 84.48 ;
      RECT  -10.93 84.25 -10.63 84.35 ;
      RECT  -7.97 83.99 -7.64 84.04 ;
      RECT  -13.73 82.61 -1.2 82.94 ;
      RECT  -12.5 85.11 -11.87 85.43 ;
      RECT  -10.93 84.04 -7.64 84.25 ;
      RECT  -5.13 84.25 -4.83 84.36 ;
      RECT  -4.74 85.35 -4.41 85.47 ;
      RECT  -10.54 84.6 -10.21 84.65 ;
      RECT  -7.97 84.25 -7.64 84.32 ;
      RECT  -12.78 84.17 -12.49 84.2 ;
      RECT  -10.54 88.58 -10.21 88.57 ;
      RECT  -12.78 89.52 -11.33 89.32 ;
      RECT  -10.54 88.82 -10.21 88.79 ;
      RECT  -4.74 88.58 -4.41 88.57 ;
      RECT  -12.78 89.32 -12.49 89.26 ;
      RECT  -3.6 88.92 -2.97 88.6 ;
      RECT  -5.82 89.24 -5.62 89.07 ;
      RECT  -5.82 88.82 -5.62 88.57 ;
      RECT  -5.13 89.67 -1.6 89.47 ;
      RECT  -10.54 89.07 -5.62 88.82 ;
      RECT  -11.62 88.57 -6.13 88.37 ;
      RECT  -11.66 89.57 -11.33 89.52 ;
      RECT  -13.65 89.43 -12.97 89.11 ;
      RECT  -6.46 88.58 -6.13 88.57 ;
      RECT  -11.66 89.32 -11.33 89.24 ;
      RECT  -13.67 87.02 -1.02 86.69 ;
      RECT  -1.94 89.77 -1.6 89.67 ;
      RECT  -10.54 88.37 -10.21 88.25 ;
      RECT  -1.94 89.47 -1.6 89.44 ;
      RECT  -11.62 89.24 -11.42 88.57 ;
      RECT  -5.82 88.57 -4.41 88.37 ;
      RECT  -6.46 88.37 -6.13 88.25 ;
      RECT  -5.86 89.57 -5.53 89.24 ;
      RECT  -10.93 89.47 -10.63 89.37 ;
      RECT  -7.97 89.73 -7.64 89.68 ;
      RECT  -13.73 91.11 -1.2 90.78 ;
      RECT  -12.5 88.61 -11.87 88.29 ;
      RECT  -10.93 89.68 -7.64 89.47 ;
      RECT  -5.13 89.47 -4.83 89.36 ;
      RECT  -4.74 88.37 -4.41 88.25 ;
      RECT  -10.54 89.12 -10.21 89.07 ;
      RECT  -7.97 89.47 -7.64 89.4 ;
      RECT  -12.78 89.55 -12.49 89.52 ;
      RECT  -10.54 93.26 -10.21 93.27 ;
      RECT  -12.78 92.32 -11.33 92.52 ;
      RECT  -10.54 93.02 -10.21 93.05 ;
      RECT  -4.74 93.26 -4.41 93.27 ;
      RECT  -12.78 92.52 -12.49 92.58 ;
      RECT  -3.6 92.92 -2.97 93.24 ;
      RECT  -5.82 92.6 -5.62 92.77 ;
      RECT  -5.82 93.02 -5.62 93.27 ;
      RECT  -5.13 92.17 -1.6 92.37 ;
      RECT  -10.54 92.77 -5.62 93.02 ;
      RECT  -11.62 93.27 -6.13 93.47 ;
      RECT  -11.66 92.27 -11.33 92.32 ;
      RECT  -13.65 92.41 -12.97 92.73 ;
      RECT  -6.46 93.26 -6.13 93.27 ;
      RECT  -11.66 92.52 -11.33 92.6 ;
      RECT  -13.67 94.82 -1.02 95.15 ;
      RECT  -1.94 92.07 -1.6 92.17 ;
      RECT  -10.54 93.47 -10.21 93.59 ;
      RECT  -1.94 92.37 -1.6 92.4 ;
      RECT  -11.62 92.6 -11.42 93.27 ;
      RECT  -5.82 93.27 -4.41 93.47 ;
      RECT  -6.46 93.47 -6.13 93.59 ;
      RECT  -5.86 92.27 -5.53 92.6 ;
      RECT  -10.93 92.37 -10.63 92.47 ;
      RECT  -7.97 92.11 -7.64 92.16 ;
      RECT  -13.73 90.73 -1.2 91.06 ;
      RECT  -12.5 93.23 -11.87 93.55 ;
      RECT  -10.93 92.16 -7.64 92.37 ;
      RECT  -5.13 92.37 -4.83 92.48 ;
      RECT  -4.74 93.47 -4.41 93.59 ;
      RECT  -10.54 92.72 -10.21 92.77 ;
      RECT  -7.97 92.37 -7.64 92.44 ;
      RECT  -12.78 92.29 -12.49 92.32 ;
      RECT  -10.54 96.7 -10.21 96.69 ;
      RECT  -12.78 97.64 -11.33 97.44 ;
      RECT  -10.54 96.94 -10.21 96.91 ;
      RECT  -4.74 96.7 -4.41 96.69 ;
      RECT  -12.78 97.44 -12.49 97.38 ;
      RECT  -3.6 97.04 -2.97 96.72 ;
      RECT  -5.82 97.36 -5.62 97.19 ;
      RECT  -5.82 96.94 -5.62 96.69 ;
      RECT  -5.13 97.79 -1.6 97.59 ;
      RECT  -10.54 97.19 -5.62 96.94 ;
      RECT  -11.62 96.69 -6.13 96.49 ;
      RECT  -11.66 97.69 -11.33 97.64 ;
      RECT  -13.65 97.55 -12.97 97.23 ;
      RECT  -6.46 96.7 -6.13 96.69 ;
      RECT  -11.66 97.44 -11.33 97.36 ;
      RECT  -13.67 95.14 -1.02 94.81 ;
      RECT  -1.94 97.89 -1.6 97.79 ;
      RECT  -10.54 96.49 -10.21 96.37 ;
      RECT  -1.94 97.59 -1.6 97.56 ;
      RECT  -11.62 97.36 -11.42 96.69 ;
      RECT  -5.82 96.69 -4.41 96.49 ;
      RECT  -6.46 96.49 -6.13 96.37 ;
      RECT  -5.86 97.69 -5.53 97.36 ;
      RECT  -10.93 97.59 -10.63 97.49 ;
      RECT  -7.97 97.85 -7.64 97.8 ;
      RECT  -13.73 99.23 -1.2 98.9 ;
      RECT  -12.5 96.73 -11.87 96.41 ;
      RECT  -10.93 97.8 -7.64 97.59 ;
      RECT  -5.13 97.59 -4.83 97.48 ;
      RECT  -4.74 96.49 -4.41 96.37 ;
      RECT  -10.54 97.24 -10.21 97.19 ;
      RECT  -7.97 97.59 -7.64 97.52 ;
      RECT  -12.78 97.67 -12.49 97.64 ;
      RECT  12.76 -7.14 13.09 -7.13 ;
      RECT  10.52 -8.08 11.97 -7.88 ;
      RECT  12.76 -7.38 13.09 -7.35 ;
      RECT  18.56 -7.14 18.89 -7.13 ;
      RECT  10.52 -7.88 10.81 -7.82 ;
      RECT  19.7 -7.48 20.33 -7.16 ;
      RECT  17.48 -7.8 17.68 -7.63 ;
      RECT  17.48 -7.38 17.68 -7.13 ;
      RECT  18.17 -8.23 21.7 -8.03 ;
      RECT  12.76 -7.63 17.68 -7.38 ;
      RECT  11.68 -7.13 17.17 -6.93 ;
      RECT  11.64 -8.13 11.97 -8.08 ;
      RECT  9.65 -7.99 10.33 -7.67 ;
      RECT  16.84 -7.14 17.17 -7.13 ;
      RECT  11.64 -7.88 11.97 -7.8 ;
      RECT  9.63 -5.58 22.28 -5.25 ;
      RECT  21.36 -8.33 21.7 -8.23 ;
      RECT  12.76 -6.93 13.09 -6.81 ;
      RECT  21.36 -8.03 21.7 -8.0 ;
      RECT  11.68 -7.8 11.88 -7.13 ;
      RECT  17.48 -7.13 18.89 -6.93 ;
      RECT  16.84 -6.93 17.17 -6.81 ;
      RECT  17.44 -8.13 17.77 -7.8 ;
      RECT  12.37 -8.03 12.67 -7.93 ;
      RECT  15.33 -8.29 15.66 -8.24 ;
      RECT  9.57 -9.67 22.1 -9.34 ;
      RECT  10.8 -7.17 11.43 -6.85 ;
      RECT  12.37 -8.24 15.66 -8.03 ;
      RECT  18.17 -8.03 18.47 -7.92 ;
      RECT  18.56 -6.93 18.89 -6.81 ;
      RECT  12.76 -7.68 13.09 -7.63 ;
      RECT  15.33 -8.03 15.66 -7.96 ;
      RECT  10.52 -8.11 10.81 -8.08 ;
      RECT  24.41 -7.14 24.74 -7.13 ;
      RECT  22.17 -8.08 23.62 -7.88 ;
      RECT  24.41 -7.38 24.74 -7.35 ;
      RECT  30.21 -7.14 30.54 -7.13 ;
      RECT  22.17 -7.88 22.46 -7.82 ;
      RECT  31.35 -7.48 31.98 -7.16 ;
      RECT  29.13 -7.8 29.33 -7.63 ;
      RECT  29.13 -7.38 29.33 -7.13 ;
      RECT  29.82 -8.23 33.35 -8.03 ;
      RECT  24.41 -7.63 29.33 -7.38 ;
      RECT  23.33 -7.13 28.82 -6.93 ;
      RECT  23.29 -8.13 23.62 -8.08 ;
      RECT  21.3 -7.99 21.98 -7.67 ;
      RECT  28.49 -7.14 28.82 -7.13 ;
      RECT  23.29 -7.88 23.62 -7.8 ;
      RECT  21.28 -5.58 33.93 -5.25 ;
      RECT  33.01 -8.33 33.35 -8.23 ;
      RECT  24.41 -6.93 24.74 -6.81 ;
      RECT  33.01 -8.03 33.35 -8.0 ;
      RECT  23.33 -7.8 23.53 -7.13 ;
      RECT  29.13 -7.13 30.54 -6.93 ;
      RECT  28.49 -6.93 28.82 -6.81 ;
      RECT  29.09 -8.13 29.42 -7.8 ;
      RECT  24.02 -8.03 24.32 -7.93 ;
      RECT  26.98 -8.29 27.31 -8.24 ;
      RECT  21.22 -9.67 33.75 -9.34 ;
      RECT  22.45 -7.17 23.08 -6.85 ;
      RECT  24.02 -8.24 27.31 -8.03 ;
      RECT  29.82 -8.03 30.12 -7.92 ;
      RECT  30.21 -6.93 30.54 -6.81 ;
      RECT  24.41 -7.68 24.74 -7.63 ;
      RECT  26.98 -8.03 27.31 -7.96 ;
      RECT  22.17 -8.11 22.46 -8.08 ;
   LAYER  m2 ;
      RECT  93.26 33.96 93.4 34.54 ;
      RECT  93.26 34.86 93.4 39.64 ;
      RECT  92.56 34.86 92.7 39.64 ;
      RECT  92.47 34.54 92.79 34.86 ;
      RECT  92.56 33.96 92.7 34.54 ;
      RECT  92.98 34.54 93.4 34.86 ;
      RECT  93.26 44.42 93.4 43.84 ;
      RECT  93.26 43.52 93.4 38.74 ;
      RECT  92.56 43.52 92.7 38.74 ;
      RECT  92.47 43.84 92.79 43.52 ;
      RECT  92.56 44.42 92.7 43.84 ;
      RECT  92.98 43.84 93.4 43.52 ;
      RECT  93.26 44.14 93.4 44.72 ;
      RECT  93.26 45.04 93.4 49.82 ;
      RECT  92.56 45.04 92.7 49.82 ;
      RECT  92.47 44.72 92.79 45.04 ;
      RECT  92.56 44.14 92.7 44.72 ;
      RECT  92.98 44.72 93.4 45.04 ;
      RECT  93.26 54.6 93.4 54.02 ;
      RECT  93.26 53.7 93.4 48.92 ;
      RECT  92.56 53.7 92.7 48.92 ;
      RECT  92.47 54.02 92.79 53.7 ;
      RECT  92.56 54.6 92.7 54.02 ;
      RECT  92.98 54.02 93.4 53.7 ;
      RECT  93.26 54.32 93.4 54.9 ;
      RECT  93.26 55.22 93.4 60.0 ;
      RECT  92.56 55.22 92.7 60.0 ;
      RECT  92.47 54.9 92.79 55.22 ;
      RECT  92.56 54.32 92.7 54.9 ;
      RECT  92.98 54.9 93.4 55.22 ;
      RECT  93.26 64.78 93.4 64.2 ;
      RECT  93.26 63.88 93.4 59.1 ;
      RECT  92.56 63.88 92.7 59.1 ;
      RECT  92.47 64.2 92.79 63.88 ;
      RECT  92.56 64.78 92.7 64.2 ;
      RECT  92.98 64.2 93.4 63.88 ;
      RECT  93.26 64.5 93.4 65.08 ;
      RECT  93.26 65.4 93.4 70.18 ;
      RECT  92.56 65.4 92.7 70.18 ;
      RECT  92.47 65.08 92.79 65.4 ;
      RECT  92.56 64.5 92.7 65.08 ;
      RECT  92.98 65.08 93.4 65.4 ;
      RECT  93.26 74.96 93.4 74.38 ;
      RECT  93.26 74.06 93.4 69.28 ;
      RECT  92.56 74.06 92.7 69.28 ;
      RECT  92.47 74.38 92.79 74.06 ;
      RECT  92.56 74.96 92.7 74.38 ;
      RECT  92.98 74.38 93.4 74.06 ;
      RECT  93.26 74.68 93.4 75.26 ;
      RECT  93.26 75.58 93.4 80.36 ;
      RECT  92.56 75.58 92.7 80.36 ;
      RECT  92.47 75.26 92.79 75.58 ;
      RECT  92.56 74.68 92.7 75.26 ;
      RECT  92.98 75.26 93.4 75.58 ;
      RECT  93.26 85.14 93.4 84.56 ;
      RECT  93.26 84.24 93.4 79.46 ;
      RECT  92.56 84.24 92.7 79.46 ;
      RECT  92.47 84.56 92.79 84.24 ;
      RECT  92.56 85.14 92.7 84.56 ;
      RECT  92.98 84.56 93.4 84.24 ;
      RECT  93.26 84.86 93.4 85.44 ;
      RECT  93.26 85.76 93.4 90.54 ;
      RECT  92.56 85.76 92.7 90.54 ;
      RECT  92.47 85.44 92.79 85.76 ;
      RECT  92.56 84.86 92.7 85.44 ;
      RECT  92.98 85.44 93.4 85.76 ;
      RECT  93.26 95.32 93.4 94.74 ;
      RECT  93.26 94.42 93.4 89.64 ;
      RECT  92.56 94.42 92.7 89.64 ;
      RECT  92.47 94.74 92.79 94.42 ;
      RECT  92.56 95.32 92.7 94.74 ;
      RECT  92.98 94.74 93.4 94.42 ;
      RECT  93.26 95.04 93.4 95.62 ;
      RECT  93.26 95.94 93.4 100.72 ;
      RECT  92.56 95.94 92.7 100.72 ;
      RECT  92.47 95.62 92.79 95.94 ;
      RECT  92.56 95.04 92.7 95.62 ;
      RECT  92.98 95.62 93.4 95.94 ;
      RECT  93.26 105.5 93.4 104.92 ;
      RECT  93.26 104.6 93.4 99.82 ;
      RECT  92.56 104.6 92.7 99.82 ;
      RECT  92.47 104.92 92.79 104.6 ;
      RECT  92.56 105.5 92.7 104.92 ;
      RECT  92.98 104.92 93.4 104.6 ;
      RECT  93.26 105.22 93.4 105.8 ;
      RECT  93.26 106.12 93.4 110.9 ;
      RECT  92.56 106.12 92.7 110.9 ;
      RECT  92.47 105.8 92.79 106.12 ;
      RECT  92.56 105.22 92.7 105.8 ;
      RECT  92.98 105.8 93.4 106.12 ;
      RECT  93.26 115.68 93.4 115.1 ;
      RECT  93.26 114.78 93.4 110.0 ;
      RECT  92.56 114.78 92.7 110.0 ;
      RECT  92.47 115.1 92.79 114.78 ;
      RECT  92.56 115.68 92.7 115.1 ;
      RECT  92.98 115.1 93.4 114.78 ;
      RECT  95.86 33.96 96.0 34.54 ;
      RECT  95.86 34.86 96.0 39.64 ;
      RECT  95.16 34.86 95.3 39.64 ;
      RECT  95.07 34.54 95.39 34.86 ;
      RECT  95.16 33.96 95.3 34.54 ;
      RECT  95.58 34.54 96.0 34.86 ;
      RECT  95.86 44.42 96.0 43.84 ;
      RECT  95.86 43.52 96.0 38.74 ;
      RECT  95.16 43.52 95.3 38.74 ;
      RECT  95.07 43.84 95.39 43.52 ;
      RECT  95.16 44.42 95.3 43.84 ;
      RECT  95.58 43.84 96.0 43.52 ;
      RECT  95.86 44.14 96.0 44.72 ;
      RECT  95.86 45.04 96.0 49.82 ;
      RECT  95.16 45.04 95.3 49.82 ;
      RECT  95.07 44.72 95.39 45.04 ;
      RECT  95.16 44.14 95.3 44.72 ;
      RECT  95.58 44.72 96.0 45.04 ;
      RECT  95.86 54.6 96.0 54.02 ;
      RECT  95.86 53.7 96.0 48.92 ;
      RECT  95.16 53.7 95.3 48.92 ;
      RECT  95.07 54.02 95.39 53.7 ;
      RECT  95.16 54.6 95.3 54.02 ;
      RECT  95.58 54.02 96.0 53.7 ;
      RECT  95.86 54.32 96.0 54.9 ;
      RECT  95.86 55.22 96.0 60.0 ;
      RECT  95.16 55.22 95.3 60.0 ;
      RECT  95.07 54.9 95.39 55.22 ;
      RECT  95.16 54.32 95.3 54.9 ;
      RECT  95.58 54.9 96.0 55.22 ;
      RECT  95.86 64.78 96.0 64.2 ;
      RECT  95.86 63.88 96.0 59.1 ;
      RECT  95.16 63.88 95.3 59.1 ;
      RECT  95.07 64.2 95.39 63.88 ;
      RECT  95.16 64.78 95.3 64.2 ;
      RECT  95.58 64.2 96.0 63.88 ;
      RECT  95.86 64.5 96.0 65.08 ;
      RECT  95.86 65.4 96.0 70.18 ;
      RECT  95.16 65.4 95.3 70.18 ;
      RECT  95.07 65.08 95.39 65.4 ;
      RECT  95.16 64.5 95.3 65.08 ;
      RECT  95.58 65.08 96.0 65.4 ;
      RECT  95.86 74.96 96.0 74.38 ;
      RECT  95.86 74.06 96.0 69.28 ;
      RECT  95.16 74.06 95.3 69.28 ;
      RECT  95.07 74.38 95.39 74.06 ;
      RECT  95.16 74.96 95.3 74.38 ;
      RECT  95.58 74.38 96.0 74.06 ;
      RECT  95.86 74.68 96.0 75.26 ;
      RECT  95.86 75.58 96.0 80.36 ;
      RECT  95.16 75.58 95.3 80.36 ;
      RECT  95.07 75.26 95.39 75.58 ;
      RECT  95.16 74.68 95.3 75.26 ;
      RECT  95.58 75.26 96.0 75.58 ;
      RECT  95.86 85.14 96.0 84.56 ;
      RECT  95.86 84.24 96.0 79.46 ;
      RECT  95.16 84.24 95.3 79.46 ;
      RECT  95.07 84.56 95.39 84.24 ;
      RECT  95.16 85.14 95.3 84.56 ;
      RECT  95.58 84.56 96.0 84.24 ;
      RECT  95.86 84.86 96.0 85.44 ;
      RECT  95.86 85.76 96.0 90.54 ;
      RECT  95.16 85.76 95.3 90.54 ;
      RECT  95.07 85.44 95.39 85.76 ;
      RECT  95.16 84.86 95.3 85.44 ;
      RECT  95.58 85.44 96.0 85.76 ;
      RECT  95.86 95.32 96.0 94.74 ;
      RECT  95.86 94.42 96.0 89.64 ;
      RECT  95.16 94.42 95.3 89.64 ;
      RECT  95.07 94.74 95.39 94.42 ;
      RECT  95.16 95.32 95.3 94.74 ;
      RECT  95.58 94.74 96.0 94.42 ;
      RECT  95.86 95.04 96.0 95.62 ;
      RECT  95.86 95.94 96.0 100.72 ;
      RECT  95.16 95.94 95.3 100.72 ;
      RECT  95.07 95.62 95.39 95.94 ;
      RECT  95.16 95.04 95.3 95.62 ;
      RECT  95.58 95.62 96.0 95.94 ;
      RECT  95.86 105.5 96.0 104.92 ;
      RECT  95.86 104.6 96.0 99.82 ;
      RECT  95.16 104.6 95.3 99.82 ;
      RECT  95.07 104.92 95.39 104.6 ;
      RECT  95.16 105.5 95.3 104.92 ;
      RECT  95.58 104.92 96.0 104.6 ;
      RECT  95.86 105.22 96.0 105.8 ;
      RECT  95.86 106.12 96.0 110.9 ;
      RECT  95.16 106.12 95.3 110.9 ;
      RECT  95.07 105.8 95.39 106.12 ;
      RECT  95.16 105.22 95.3 105.8 ;
      RECT  95.58 105.8 96.0 106.12 ;
      RECT  95.86 115.68 96.0 115.1 ;
      RECT  95.86 114.78 96.0 110.0 ;
      RECT  95.16 114.78 95.3 110.0 ;
      RECT  95.07 115.1 95.39 114.78 ;
      RECT  95.16 115.68 95.3 115.1 ;
      RECT  95.58 115.1 96.0 114.78 ;
      RECT  92.47 34.1 92.79 115.54 ;
      RECT  92.98 34.1 93.4 115.54 ;
      RECT  95.07 34.1 95.39 115.54 ;
      RECT  95.58 34.1 96.0 115.54 ;
      RECT  90.66 23.78 90.8 24.36 ;
      RECT  90.66 24.68 90.8 29.46 ;
      RECT  89.96 24.68 90.1 29.46 ;
      RECT  89.87 24.36 90.19 24.68 ;
      RECT  89.96 23.78 90.1 24.36 ;
      RECT  90.38 24.36 90.8 24.68 ;
      RECT  90.66 34.24 90.8 33.66 ;
      RECT  90.66 33.34 90.8 28.56 ;
      RECT  89.96 33.34 90.1 28.56 ;
      RECT  89.87 33.66 90.19 33.34 ;
      RECT  89.96 34.24 90.1 33.66 ;
      RECT  90.38 33.66 90.8 33.34 ;
      RECT  90.66 33.96 90.8 34.54 ;
      RECT  90.66 34.86 90.8 39.64 ;
      RECT  89.96 34.86 90.1 39.64 ;
      RECT  89.87 34.54 90.19 34.86 ;
      RECT  89.96 33.96 90.1 34.54 ;
      RECT  90.38 34.54 90.8 34.86 ;
      RECT  90.66 44.42 90.8 43.84 ;
      RECT  90.66 43.52 90.8 38.74 ;
      RECT  89.96 43.52 90.1 38.74 ;
      RECT  89.87 43.84 90.19 43.52 ;
      RECT  89.96 44.42 90.1 43.84 ;
      RECT  90.38 43.84 90.8 43.52 ;
      RECT  90.66 44.14 90.8 44.72 ;
      RECT  90.66 45.04 90.8 49.82 ;
      RECT  89.96 45.04 90.1 49.82 ;
      RECT  89.87 44.72 90.19 45.04 ;
      RECT  89.96 44.14 90.1 44.72 ;
      RECT  90.38 44.72 90.8 45.04 ;
      RECT  90.66 54.6 90.8 54.02 ;
      RECT  90.66 53.7 90.8 48.92 ;
      RECT  89.96 53.7 90.1 48.92 ;
      RECT  89.87 54.02 90.19 53.7 ;
      RECT  89.96 54.6 90.1 54.02 ;
      RECT  90.38 54.02 90.8 53.7 ;
      RECT  90.66 54.32 90.8 54.9 ;
      RECT  90.66 55.22 90.8 60.0 ;
      RECT  89.96 55.22 90.1 60.0 ;
      RECT  89.87 54.9 90.19 55.22 ;
      RECT  89.96 54.32 90.1 54.9 ;
      RECT  90.38 54.9 90.8 55.22 ;
      RECT  90.66 64.78 90.8 64.2 ;
      RECT  90.66 63.88 90.8 59.1 ;
      RECT  89.96 63.88 90.1 59.1 ;
      RECT  89.87 64.2 90.19 63.88 ;
      RECT  89.96 64.78 90.1 64.2 ;
      RECT  90.38 64.2 90.8 63.88 ;
      RECT  90.66 64.5 90.8 65.08 ;
      RECT  90.66 65.4 90.8 70.18 ;
      RECT  89.96 65.4 90.1 70.18 ;
      RECT  89.87 65.08 90.19 65.4 ;
      RECT  89.96 64.5 90.1 65.08 ;
      RECT  90.38 65.08 90.8 65.4 ;
      RECT  90.66 74.96 90.8 74.38 ;
      RECT  90.66 74.06 90.8 69.28 ;
      RECT  89.96 74.06 90.1 69.28 ;
      RECT  89.87 74.38 90.19 74.06 ;
      RECT  89.96 74.96 90.1 74.38 ;
      RECT  90.38 74.38 90.8 74.06 ;
      RECT  90.66 74.68 90.8 75.26 ;
      RECT  90.66 75.58 90.8 80.36 ;
      RECT  89.96 75.58 90.1 80.36 ;
      RECT  89.87 75.26 90.19 75.58 ;
      RECT  89.96 74.68 90.1 75.26 ;
      RECT  90.38 75.26 90.8 75.58 ;
      RECT  90.66 85.14 90.8 84.56 ;
      RECT  90.66 84.24 90.8 79.46 ;
      RECT  89.96 84.24 90.1 79.46 ;
      RECT  89.87 84.56 90.19 84.24 ;
      RECT  89.96 85.14 90.1 84.56 ;
      RECT  90.38 84.56 90.8 84.24 ;
      RECT  90.66 84.86 90.8 85.44 ;
      RECT  90.66 85.76 90.8 90.54 ;
      RECT  89.96 85.76 90.1 90.54 ;
      RECT  89.87 85.44 90.19 85.76 ;
      RECT  89.96 84.86 90.1 85.44 ;
      RECT  90.38 85.44 90.8 85.76 ;
      RECT  90.66 95.32 90.8 94.74 ;
      RECT  90.66 94.42 90.8 89.64 ;
      RECT  89.96 94.42 90.1 89.64 ;
      RECT  89.87 94.74 90.19 94.42 ;
      RECT  89.96 95.32 90.1 94.74 ;
      RECT  90.38 94.74 90.8 94.42 ;
      RECT  90.66 95.04 90.8 95.62 ;
      RECT  90.66 95.94 90.8 100.72 ;
      RECT  89.96 95.94 90.1 100.72 ;
      RECT  89.87 95.62 90.19 95.94 ;
      RECT  89.96 95.04 90.1 95.62 ;
      RECT  90.38 95.62 90.8 95.94 ;
      RECT  90.66 105.5 90.8 104.92 ;
      RECT  90.66 104.6 90.8 99.82 ;
      RECT  89.96 104.6 90.1 99.82 ;
      RECT  89.87 104.92 90.19 104.6 ;
      RECT  89.96 105.5 90.1 104.92 ;
      RECT  90.38 104.92 90.8 104.6 ;
      RECT  90.66 105.22 90.8 105.8 ;
      RECT  90.66 106.12 90.8 110.9 ;
      RECT  89.96 106.12 90.1 110.9 ;
      RECT  89.87 105.8 90.19 106.12 ;
      RECT  89.96 105.22 90.1 105.8 ;
      RECT  90.38 105.8 90.8 106.12 ;
      RECT  90.66 115.68 90.8 115.1 ;
      RECT  90.66 114.78 90.8 110.0 ;
      RECT  89.96 114.78 90.1 110.0 ;
      RECT  89.87 115.1 90.19 114.78 ;
      RECT  89.96 115.68 90.1 115.1 ;
      RECT  90.38 115.1 90.8 114.78 ;
      RECT  90.66 115.4 90.8 115.98 ;
      RECT  90.66 116.3 90.8 121.08 ;
      RECT  89.96 116.3 90.1 121.08 ;
      RECT  89.87 115.98 90.19 116.3 ;
      RECT  89.96 115.4 90.1 115.98 ;
      RECT  90.38 115.98 90.8 116.3 ;
      RECT  89.87 23.92 90.19 120.63 ;
      RECT  90.38 23.92 90.8 120.63 ;
      RECT  93.26 34.24 93.4 33.66 ;
      RECT  93.26 33.34 93.4 28.56 ;
      RECT  92.56 33.34 92.7 28.56 ;
      RECT  92.47 33.66 92.79 33.34 ;
      RECT  92.56 34.24 92.7 33.66 ;
      RECT  92.98 33.66 93.4 33.34 ;
      RECT  95.86 34.24 96.0 33.66 ;
      RECT  95.86 33.34 96.0 28.56 ;
      RECT  95.16 33.34 95.3 28.56 ;
      RECT  95.07 33.66 95.39 33.34 ;
      RECT  95.16 34.24 95.3 33.66 ;
      RECT  95.58 33.66 96.0 33.34 ;
      RECT  92.47 34.1 92.79 29.01 ;
      RECT  92.98 34.1 93.4 29.01 ;
      RECT  95.07 34.1 95.39 29.01 ;
      RECT  95.58 34.1 96.0 29.01 ;
      RECT  93.26 23.78 93.4 24.36 ;
      RECT  93.26 24.68 93.4 29.46 ;
      RECT  92.56 24.68 92.7 29.46 ;
      RECT  92.47 24.36 92.79 24.68 ;
      RECT  92.56 23.78 92.7 24.36 ;
      RECT  92.98 24.36 93.4 24.68 ;
      RECT  95.86 23.78 96.0 24.36 ;
      RECT  95.86 24.68 96.0 29.46 ;
      RECT  95.16 24.68 95.3 29.46 ;
      RECT  95.07 24.36 95.39 24.68 ;
      RECT  95.16 23.78 95.3 24.36 ;
      RECT  95.58 24.36 96.0 24.68 ;
      RECT  92.47 23.92 92.79 29.01 ;
      RECT  92.98 23.92 93.4 29.01 ;
      RECT  95.07 23.92 95.39 29.01 ;
      RECT  95.58 23.92 96.0 29.01 ;
      RECT  93.26 115.4 93.4 115.98 ;
      RECT  93.26 116.3 93.4 121.08 ;
      RECT  92.56 116.3 92.7 121.08 ;
      RECT  92.47 115.98 92.79 116.3 ;
      RECT  92.56 115.4 92.7 115.98 ;
      RECT  92.98 115.98 93.4 116.3 ;
      RECT  95.86 115.4 96.0 115.98 ;
      RECT  95.86 116.3 96.0 121.08 ;
      RECT  95.16 116.3 95.3 121.08 ;
      RECT  95.07 115.98 95.39 116.3 ;
      RECT  95.16 115.4 95.3 115.98 ;
      RECT  95.58 115.98 96.0 116.3 ;
      RECT  92.47 115.54 92.79 120.63 ;
      RECT  92.98 115.54 93.4 120.63 ;
      RECT  95.07 115.54 95.39 120.63 ;
      RECT  95.58 115.54 96.0 120.63 ;
      RECT  88.06 23.78 88.2 24.36 ;
      RECT  88.06 24.68 88.2 29.46 ;
      RECT  87.36 24.68 87.5 29.46 ;
      RECT  87.27 24.36 87.59 24.68 ;
      RECT  87.36 23.78 87.5 24.36 ;
      RECT  87.78 24.36 88.2 24.68 ;
      RECT  88.06 34.24 88.2 33.66 ;
      RECT  88.06 33.34 88.2 28.56 ;
      RECT  87.36 33.34 87.5 28.56 ;
      RECT  87.27 33.66 87.59 33.34 ;
      RECT  87.36 34.24 87.5 33.66 ;
      RECT  87.78 33.66 88.2 33.34 ;
      RECT  88.06 33.96 88.2 34.54 ;
      RECT  88.06 34.86 88.2 39.64 ;
      RECT  87.36 34.86 87.5 39.64 ;
      RECT  87.27 34.54 87.59 34.86 ;
      RECT  87.36 33.96 87.5 34.54 ;
      RECT  87.78 34.54 88.2 34.86 ;
      RECT  88.06 44.42 88.2 43.84 ;
      RECT  88.06 43.52 88.2 38.74 ;
      RECT  87.36 43.52 87.5 38.74 ;
      RECT  87.27 43.84 87.59 43.52 ;
      RECT  87.36 44.42 87.5 43.84 ;
      RECT  87.78 43.84 88.2 43.52 ;
      RECT  88.06 44.14 88.2 44.72 ;
      RECT  88.06 45.04 88.2 49.82 ;
      RECT  87.36 45.04 87.5 49.82 ;
      RECT  87.27 44.72 87.59 45.04 ;
      RECT  87.36 44.14 87.5 44.72 ;
      RECT  87.78 44.72 88.2 45.04 ;
      RECT  88.06 54.6 88.2 54.02 ;
      RECT  88.06 53.7 88.2 48.92 ;
      RECT  87.36 53.7 87.5 48.92 ;
      RECT  87.27 54.02 87.59 53.7 ;
      RECT  87.36 54.6 87.5 54.02 ;
      RECT  87.78 54.02 88.2 53.7 ;
      RECT  88.06 54.32 88.2 54.9 ;
      RECT  88.06 55.22 88.2 60.0 ;
      RECT  87.36 55.22 87.5 60.0 ;
      RECT  87.27 54.9 87.59 55.22 ;
      RECT  87.36 54.32 87.5 54.9 ;
      RECT  87.78 54.9 88.2 55.22 ;
      RECT  88.06 64.78 88.2 64.2 ;
      RECT  88.06 63.88 88.2 59.1 ;
      RECT  87.36 63.88 87.5 59.1 ;
      RECT  87.27 64.2 87.59 63.88 ;
      RECT  87.36 64.78 87.5 64.2 ;
      RECT  87.78 64.2 88.2 63.88 ;
      RECT  88.06 64.5 88.2 65.08 ;
      RECT  88.06 65.4 88.2 70.18 ;
      RECT  87.36 65.4 87.5 70.18 ;
      RECT  87.27 65.08 87.59 65.4 ;
      RECT  87.36 64.5 87.5 65.08 ;
      RECT  87.78 65.08 88.2 65.4 ;
      RECT  88.06 74.96 88.2 74.38 ;
      RECT  88.06 74.06 88.2 69.28 ;
      RECT  87.36 74.06 87.5 69.28 ;
      RECT  87.27 74.38 87.59 74.06 ;
      RECT  87.36 74.96 87.5 74.38 ;
      RECT  87.78 74.38 88.2 74.06 ;
      RECT  88.06 74.68 88.2 75.26 ;
      RECT  88.06 75.58 88.2 80.36 ;
      RECT  87.36 75.58 87.5 80.36 ;
      RECT  87.27 75.26 87.59 75.58 ;
      RECT  87.36 74.68 87.5 75.26 ;
      RECT  87.78 75.26 88.2 75.58 ;
      RECT  88.06 85.14 88.2 84.56 ;
      RECT  88.06 84.24 88.2 79.46 ;
      RECT  87.36 84.24 87.5 79.46 ;
      RECT  87.27 84.56 87.59 84.24 ;
      RECT  87.36 85.14 87.5 84.56 ;
      RECT  87.78 84.56 88.2 84.24 ;
      RECT  88.06 84.86 88.2 85.44 ;
      RECT  88.06 85.76 88.2 90.54 ;
      RECT  87.36 85.76 87.5 90.54 ;
      RECT  87.27 85.44 87.59 85.76 ;
      RECT  87.36 84.86 87.5 85.44 ;
      RECT  87.78 85.44 88.2 85.76 ;
      RECT  88.06 95.32 88.2 94.74 ;
      RECT  88.06 94.42 88.2 89.64 ;
      RECT  87.36 94.42 87.5 89.64 ;
      RECT  87.27 94.74 87.59 94.42 ;
      RECT  87.36 95.32 87.5 94.74 ;
      RECT  87.78 94.74 88.2 94.42 ;
      RECT  88.06 95.04 88.2 95.62 ;
      RECT  88.06 95.94 88.2 100.72 ;
      RECT  87.36 95.94 87.5 100.72 ;
      RECT  87.27 95.62 87.59 95.94 ;
      RECT  87.36 95.04 87.5 95.62 ;
      RECT  87.78 95.62 88.2 95.94 ;
      RECT  88.06 105.5 88.2 104.92 ;
      RECT  88.06 104.6 88.2 99.82 ;
      RECT  87.36 104.6 87.5 99.82 ;
      RECT  87.27 104.92 87.59 104.6 ;
      RECT  87.36 105.5 87.5 104.92 ;
      RECT  87.78 104.92 88.2 104.6 ;
      RECT  88.06 105.22 88.2 105.8 ;
      RECT  88.06 106.12 88.2 110.9 ;
      RECT  87.36 106.12 87.5 110.9 ;
      RECT  87.27 105.8 87.59 106.12 ;
      RECT  87.36 105.22 87.5 105.8 ;
      RECT  87.78 105.8 88.2 106.12 ;
      RECT  88.06 115.68 88.2 115.1 ;
      RECT  88.06 114.78 88.2 110.0 ;
      RECT  87.36 114.78 87.5 110.0 ;
      RECT  87.27 115.1 87.59 114.78 ;
      RECT  87.36 115.68 87.5 115.1 ;
      RECT  87.78 115.1 88.2 114.78 ;
      RECT  88.06 115.4 88.2 115.98 ;
      RECT  88.06 116.3 88.2 121.08 ;
      RECT  87.36 116.3 87.5 121.08 ;
      RECT  87.27 115.98 87.59 116.3 ;
      RECT  87.36 115.4 87.5 115.98 ;
      RECT  87.78 115.98 88.2 116.3 ;
      RECT  87.27 23.92 87.59 120.63 ;
      RECT  87.78 23.92 88.2 120.63 ;
      RECT  98.46 23.78 98.6 24.36 ;
      RECT  98.46 24.68 98.6 29.46 ;
      RECT  97.76 24.68 97.9 29.46 ;
      RECT  97.67 24.36 97.99 24.68 ;
      RECT  97.76 23.78 97.9 24.36 ;
      RECT  98.18 24.36 98.6 24.68 ;
      RECT  98.46 34.24 98.6 33.66 ;
      RECT  98.46 33.34 98.6 28.56 ;
      RECT  97.76 33.34 97.9 28.56 ;
      RECT  97.67 33.66 97.99 33.34 ;
      RECT  97.76 34.24 97.9 33.66 ;
      RECT  98.18 33.66 98.6 33.34 ;
      RECT  98.46 33.96 98.6 34.54 ;
      RECT  98.46 34.86 98.6 39.64 ;
      RECT  97.76 34.86 97.9 39.64 ;
      RECT  97.67 34.54 97.99 34.86 ;
      RECT  97.76 33.96 97.9 34.54 ;
      RECT  98.18 34.54 98.6 34.86 ;
      RECT  98.46 44.42 98.6 43.84 ;
      RECT  98.46 43.52 98.6 38.74 ;
      RECT  97.76 43.52 97.9 38.74 ;
      RECT  97.67 43.84 97.99 43.52 ;
      RECT  97.76 44.42 97.9 43.84 ;
      RECT  98.18 43.84 98.6 43.52 ;
      RECT  98.46 44.14 98.6 44.72 ;
      RECT  98.46 45.04 98.6 49.82 ;
      RECT  97.76 45.04 97.9 49.82 ;
      RECT  97.67 44.72 97.99 45.04 ;
      RECT  97.76 44.14 97.9 44.72 ;
      RECT  98.18 44.72 98.6 45.04 ;
      RECT  98.46 54.6 98.6 54.02 ;
      RECT  98.46 53.7 98.6 48.92 ;
      RECT  97.76 53.7 97.9 48.92 ;
      RECT  97.67 54.02 97.99 53.7 ;
      RECT  97.76 54.6 97.9 54.02 ;
      RECT  98.18 54.02 98.6 53.7 ;
      RECT  98.46 54.32 98.6 54.9 ;
      RECT  98.46 55.22 98.6 60.0 ;
      RECT  97.76 55.22 97.9 60.0 ;
      RECT  97.67 54.9 97.99 55.22 ;
      RECT  97.76 54.32 97.9 54.9 ;
      RECT  98.18 54.9 98.6 55.22 ;
      RECT  98.46 64.78 98.6 64.2 ;
      RECT  98.46 63.88 98.6 59.1 ;
      RECT  97.76 63.88 97.9 59.1 ;
      RECT  97.67 64.2 97.99 63.88 ;
      RECT  97.76 64.78 97.9 64.2 ;
      RECT  98.18 64.2 98.6 63.88 ;
      RECT  98.46 64.5 98.6 65.08 ;
      RECT  98.46 65.4 98.6 70.18 ;
      RECT  97.76 65.4 97.9 70.18 ;
      RECT  97.67 65.08 97.99 65.4 ;
      RECT  97.76 64.5 97.9 65.08 ;
      RECT  98.18 65.08 98.6 65.4 ;
      RECT  98.46 74.96 98.6 74.38 ;
      RECT  98.46 74.06 98.6 69.28 ;
      RECT  97.76 74.06 97.9 69.28 ;
      RECT  97.67 74.38 97.99 74.06 ;
      RECT  97.76 74.96 97.9 74.38 ;
      RECT  98.18 74.38 98.6 74.06 ;
      RECT  98.46 74.68 98.6 75.26 ;
      RECT  98.46 75.58 98.6 80.36 ;
      RECT  97.76 75.58 97.9 80.36 ;
      RECT  97.67 75.26 97.99 75.58 ;
      RECT  97.76 74.68 97.9 75.26 ;
      RECT  98.18 75.26 98.6 75.58 ;
      RECT  98.46 85.14 98.6 84.56 ;
      RECT  98.46 84.24 98.6 79.46 ;
      RECT  97.76 84.24 97.9 79.46 ;
      RECT  97.67 84.56 97.99 84.24 ;
      RECT  97.76 85.14 97.9 84.56 ;
      RECT  98.18 84.56 98.6 84.24 ;
      RECT  98.46 84.86 98.6 85.44 ;
      RECT  98.46 85.76 98.6 90.54 ;
      RECT  97.76 85.76 97.9 90.54 ;
      RECT  97.67 85.44 97.99 85.76 ;
      RECT  97.76 84.86 97.9 85.44 ;
      RECT  98.18 85.44 98.6 85.76 ;
      RECT  98.46 95.32 98.6 94.74 ;
      RECT  98.46 94.42 98.6 89.64 ;
      RECT  97.76 94.42 97.9 89.64 ;
      RECT  97.67 94.74 97.99 94.42 ;
      RECT  97.76 95.32 97.9 94.74 ;
      RECT  98.18 94.74 98.6 94.42 ;
      RECT  98.46 95.04 98.6 95.62 ;
      RECT  98.46 95.94 98.6 100.72 ;
      RECT  97.76 95.94 97.9 100.72 ;
      RECT  97.67 95.62 97.99 95.94 ;
      RECT  97.76 95.04 97.9 95.62 ;
      RECT  98.18 95.62 98.6 95.94 ;
      RECT  98.46 105.5 98.6 104.92 ;
      RECT  98.46 104.6 98.6 99.82 ;
      RECT  97.76 104.6 97.9 99.82 ;
      RECT  97.67 104.92 97.99 104.6 ;
      RECT  97.76 105.5 97.9 104.92 ;
      RECT  98.18 104.92 98.6 104.6 ;
      RECT  98.46 105.22 98.6 105.8 ;
      RECT  98.46 106.12 98.6 110.9 ;
      RECT  97.76 106.12 97.9 110.9 ;
      RECT  97.67 105.8 97.99 106.12 ;
      RECT  97.76 105.22 97.9 105.8 ;
      RECT  98.18 105.8 98.6 106.12 ;
      RECT  98.46 115.68 98.6 115.1 ;
      RECT  98.46 114.78 98.6 110.0 ;
      RECT  97.76 114.78 97.9 110.0 ;
      RECT  97.67 115.1 97.99 114.78 ;
      RECT  97.76 115.68 97.9 115.1 ;
      RECT  98.18 115.1 98.6 114.78 ;
      RECT  98.46 115.4 98.6 115.98 ;
      RECT  98.46 116.3 98.6 121.08 ;
      RECT  97.76 116.3 97.9 121.08 ;
      RECT  97.67 115.98 97.99 116.3 ;
      RECT  97.76 115.4 97.9 115.98 ;
      RECT  98.18 115.98 98.6 116.3 ;
      RECT  97.67 23.92 97.99 120.63 ;
      RECT  98.18 23.92 98.6 120.63 ;
      RECT  89.87 23.92 90.19 120.63 ;
      RECT  90.38 23.92 90.8 120.63 ;
      RECT  92.47 23.92 92.79 120.63 ;
      RECT  92.98 23.92 93.4 120.63 ;
      RECT  95.07 23.92 95.39 120.63 ;
      RECT  95.58 23.92 96.0 120.63 ;
      RECT  89.45 14.29 89.59 22.39 ;
      RECT  91.03 14.29 91.17 22.39 ;
      RECT  92.05 14.29 92.19 22.39 ;
      RECT  93.63 14.29 93.77 22.39 ;
      RECT  94.65 14.29 94.79 22.39 ;
      RECT  96.23 14.29 96.37 22.39 ;
      RECT  89.45 14.29 89.59 22.39 ;
      RECT  91.03 14.29 91.17 22.39 ;
      RECT  92.05 14.29 92.19 22.39 ;
      RECT  93.63 14.29 93.77 22.39 ;
      RECT  94.65 14.29 94.79 22.39 ;
      RECT  96.23 14.29 96.37 22.39 ;
      RECT  91.32 8.18 91.65 13.22 ;
      RECT  96.9 8.18 97.23 13.22 ;
      RECT  92.96 8.18 93.29 13.22 ;
      RECT  93.92 8.18 94.25 13.22 ;
      RECT  99.5 8.18 99.83 13.22 ;
      RECT  95.56 8.18 95.89 13.22 ;
      RECT  89.45 22.39 89.59 14.29 ;
      RECT  91.03 22.39 91.17 14.29 ;
      RECT  92.05 22.39 92.19 14.29 ;
      RECT  93.63 22.39 93.77 14.29 ;
      RECT  94.65 22.39 94.79 14.29 ;
      RECT  96.23 22.39 96.37 14.29 ;
      RECT  2.69 36.38 3.01 36.7 ;
      RECT  3.2 41.68 3.52 42.0 ;
      RECT  2.69 66.92 3.01 67.24 ;
      RECT  3.2 72.22 3.52 72.54 ;
      RECT  0.09 34.1 0.23 85.0 ;
      RECT  0.6 34.1 0.74 85.0 ;
      RECT  1.11 34.1 1.25 85.0 ;
      RECT  1.62 34.1 1.76 85.0 ;
      RECT  70.46 34.1 70.6 115.54 ;
      RECT  0.09 34.1 0.23 85.0 ;
      RECT  0.6 34.1 0.74 85.0 ;
      RECT  1.11 34.1 1.25 85.0 ;
      RECT  1.62 34.1 1.76 85.0 ;
      RECT  66.26 32.56 66.4 32.7 ;
      RECT  0.09 34.1 0.23 85.0 ;
      RECT  0.6 34.1 0.74 85.0 ;
      RECT  1.11 34.1 1.25 85.0 ;
      RECT  1.62 34.1 1.76 85.0 ;
      RECT  81.64 0.0 81.78 23.92 ;
      RECT  83.0 0.0 83.14 23.92 ;
      RECT  82.32 0.0 82.46 23.92 ;
      RECT  83.68 0.0 83.82 23.92 ;
      RECT  -102.14 -7.17 -101.8 -6.85 ;
      RECT  -93.24 -7.48 -92.92 -7.16 ;
      RECT  -102.92 -7.99 -102.61 -7.67 ;
      RECT  -102.14 -7.17 -101.8 -6.85 ;
      RECT  -70.5 -8.68 -70.36 -8.54 ;
      RECT  -79.92 -6.61 -79.78 -6.47 ;
      RECT  -102.92 -7.99 -102.61 -7.67 ;
      RECT  -102.14 -3.67 -101.8 -3.99 ;
      RECT  -93.24 -3.36 -92.92 -3.68 ;
      RECT  -102.92 -2.85 -102.61 -3.17 ;
      RECT  -102.14 -3.67 -101.8 -3.99 ;
      RECT  -70.5 -2.16 -70.36 -2.3 ;
      RECT  -79.92 -4.23 -79.78 -4.37 ;
      RECT  -102.92 -2.85 -102.61 -3.17 ;
      RECT  -102.14 -7.17 -101.8 -6.85 ;
      RECT  -102.14 -3.99 -101.8 -3.67 ;
      RECT  -70.5 -8.68 -70.36 -8.54 ;
      RECT  -79.92 -6.61 -79.78 -6.47 ;
      RECT  -70.5 -2.3 -70.36 -2.16 ;
      RECT  -79.92 -4.37 -79.78 -4.23 ;
      RECT  -102.92 -9.48 -102.78 -1.36 ;
      RECT  -63.2 23.92 -63.34 27.03 ;
      RECT  -97.47 23.92 -97.61 78.55 ;
      RECT  -102.14 -7.17 -101.8 -6.85 ;
      RECT  -102.14 -3.99 -101.8 -3.67 ;
      RECT  -57.65 -7.63 -57.51 -7.49 ;
      RECT  -63.34 23.92 -63.2 27.03 ;
      RECT  -40.52 21.01 -1.02 21.15 ;
      RECT  -33.12 8.57 -1.02 8.71 ;
      RECT  -33.93 12.89 -1.02 13.03 ;
      RECT  -29.09 4.79 -1.02 4.93 ;
      RECT  -15.29 -7.68 -1.02 -7.54 ;
      RECT  -12.5 85.11 -12.16 85.43 ;
      RECT  -3.6 84.8 -3.28 85.12 ;
      RECT  -13.28 84.29 -12.97 84.61 ;
      RECT  -12.5 88.61 -12.16 88.29 ;
      RECT  -3.6 88.92 -3.28 88.6 ;
      RECT  -13.28 89.43 -12.97 89.11 ;
      RECT  -12.5 93.23 -12.16 93.55 ;
      RECT  -3.6 92.92 -3.28 93.24 ;
      RECT  -13.28 92.41 -12.97 92.73 ;
      RECT  -12.5 96.73 -12.16 96.41 ;
      RECT  -3.6 97.04 -3.28 96.72 ;
      RECT  -13.28 97.55 -12.97 97.23 ;
      RECT  -12.5 85.11 -12.16 85.43 ;
      RECT  -12.5 88.29 -12.16 88.61 ;
      RECT  -12.5 93.23 -12.16 93.55 ;
      RECT  -12.5 96.41 -12.16 96.73 ;
      RECT  -3.6 84.8 -3.28 85.12 ;
      RECT  -3.6 88.6 -3.28 88.92 ;
      RECT  -3.6 92.92 -3.28 93.24 ;
      RECT  -3.6 96.72 -3.28 97.04 ;
      RECT  10.8 -7.17 11.14 -6.85 ;
      RECT  19.7 -7.48 20.02 -7.16 ;
      RECT  10.02 -7.99 10.33 -7.67 ;
      RECT  22.45 -7.17 22.79 -6.85 ;
      RECT  31.35 -7.48 31.67 -7.16 ;
      RECT  21.67 -7.99 21.98 -7.67 ;
      RECT  10.8 -7.17 11.14 -6.85 ;
      RECT  22.45 -7.17 22.79 -6.85 ;
      RECT  19.7 -7.48 20.02 -7.16 ;
      RECT  31.35 -7.48 31.67 -7.16 ;
   LAYER  m3 ;
      RECT  90.13 28.82 90.49 29.19 ;
      RECT  90.13 120.44 90.49 120.81 ;
      RECT  90.13 23.74 90.49 24.11 ;
      RECT  90.13 115.36 90.49 115.73 ;
      RECT  97.92 28.83 98.3 29.2 ;
      RECT  97.92 100.08 98.3 100.45 ;
      RECT  97.92 120.44 98.3 120.81 ;
      RECT  87.52 49.19 87.9 49.56 ;
      RECT  92.72 120.44 93.1 120.81 ;
      RECT  97.92 28.82 98.3 29.19 ;
      RECT  87.52 100.09 87.9 100.46 ;
      RECT  87.52 49.18 87.9 49.55 ;
      RECT  97.92 39.0 98.3 39.37 ;
      RECT  95.32 120.44 95.7 120.81 ;
      RECT  87.52 79.72 87.9 80.09 ;
      RECT  87.52 100.08 87.9 100.45 ;
      RECT  87.52 89.9 87.9 90.27 ;
      RECT  87.52 120.44 87.9 120.81 ;
      RECT  87.52 39.0 87.9 39.37 ;
      RECT  87.52 79.73 87.9 80.1 ;
      RECT  87.52 28.82 87.9 29.19 ;
      RECT  95.32 28.82 95.7 29.19 ;
      RECT  90.13 28.82 90.49 29.19 ;
      RECT  97.92 49.19 98.3 49.56 ;
      RECT  87.52 59.36 87.9 59.73 ;
      RECT  97.92 59.37 98.3 59.74 ;
      RECT  97.92 110.26 98.3 110.63 ;
      RECT  87.52 110.27 87.9 110.64 ;
      RECT  87.52 39.01 87.9 39.38 ;
      RECT  97.92 69.55 98.3 69.92 ;
      RECT  87.52 69.55 87.9 69.92 ;
      RECT  87.52 89.91 87.9 90.28 ;
      RECT  97.92 100.09 98.3 100.46 ;
      RECT  87.52 69.54 87.9 69.91 ;
      RECT  92.72 28.82 93.1 29.19 ;
      RECT  97.92 79.73 98.3 80.1 ;
      RECT  97.92 89.9 98.3 90.27 ;
      RECT  87.52 59.37 87.9 59.74 ;
      RECT  97.92 69.54 98.3 69.91 ;
      RECT  97.92 79.72 98.3 80.09 ;
      RECT  97.92 59.36 98.3 59.73 ;
      RECT  97.92 89.91 98.3 90.28 ;
      RECT  97.92 110.27 98.3 110.64 ;
      RECT  87.52 110.26 87.9 110.63 ;
      RECT  90.13 120.44 90.49 120.81 ;
      RECT  97.92 49.18 98.3 49.55 ;
      RECT  97.92 39.01 98.3 39.38 ;
      RECT  87.52 28.83 87.9 29.2 ;
      RECT  97.92 64.46 98.3 64.83 ;
      RECT  97.92 74.63 98.3 75.0 ;
      RECT  97.92 33.92 98.3 34.29 ;
      RECT  87.52 54.28 87.9 54.65 ;
      RECT  87.52 94.99 87.9 95.36 ;
      RECT  97.92 64.45 98.3 64.82 ;
      RECT  87.52 95.0 87.9 95.37 ;
      RECT  97.92 44.09 98.3 44.46 ;
      RECT  99.92 24.88 100.28 25.26 ;
      RECT  87.52 115.35 87.9 115.72 ;
      RECT  99.92 116.5 100.28 116.88 ;
      RECT  97.92 54.28 98.3 54.65 ;
      RECT  97.92 84.82 98.3 85.19 ;
      RECT  92.72 23.74 93.1 24.11 ;
      RECT  85.54 24.88 85.9 25.26 ;
      RECT  87.52 74.63 87.9 75.0 ;
      RECT  87.52 105.18 87.9 105.55 ;
      RECT  87.52 44.1 87.9 44.47 ;
      RECT  97.92 105.18 98.3 105.55 ;
      RECT  87.52 64.45 87.9 64.82 ;
      RECT  90.13 23.74 90.49 24.11 ;
      RECT  97.92 105.17 98.3 105.54 ;
      RECT  97.92 74.64 98.3 75.01 ;
      RECT  87.52 84.81 87.9 85.18 ;
      RECT  95.32 115.36 95.7 115.73 ;
      RECT  97.92 95.0 98.3 95.37 ;
      RECT  97.92 115.36 98.3 115.73 ;
      RECT  95.32 23.74 95.7 24.11 ;
      RECT  87.52 33.91 87.9 34.28 ;
      RECT  97.92 44.1 98.3 44.47 ;
      RECT  97.92 33.91 98.3 34.28 ;
      RECT  87.52 64.46 87.9 64.83 ;
      RECT  87.52 23.74 87.9 24.11 ;
      RECT  97.92 54.27 98.3 54.64 ;
      RECT  90.13 115.36 90.49 115.73 ;
      RECT  97.92 84.81 98.3 85.18 ;
      RECT  87.52 44.09 87.9 44.46 ;
      RECT  87.52 74.64 87.9 75.01 ;
      RECT  87.52 115.36 87.9 115.73 ;
      RECT  87.52 105.17 87.9 105.54 ;
      RECT  97.92 115.35 98.3 115.72 ;
      RECT  87.52 54.27 87.9 54.64 ;
      RECT  92.72 115.36 93.1 115.73 ;
      RECT  97.92 94.99 98.3 95.36 ;
      RECT  85.54 116.5 85.9 116.88 ;
      RECT  87.52 84.82 87.9 85.19 ;
      RECT  87.52 33.92 87.9 34.29 ;
      RECT  97.92 23.74 98.3 24.11 ;
      RECT  94.54 19.91 94.91 20.29 ;
      RECT  97.14 19.91 97.51 20.29 ;
      RECT  99.74 19.91 100.11 20.29 ;
      RECT  97.14 19.91 97.51 20.29 ;
      RECT  99.74 19.91 100.11 20.29 ;
      RECT  94.54 19.91 94.91 20.29 ;
      RECT  96.76 12.57 97.13 12.94 ;
      RECT  94.16 12.57 94.53 12.94 ;
      RECT  94.16 8.2 94.53 8.57 ;
      RECT  96.76 8.2 97.13 8.57 ;
      RECT  98.72 6.98 99.08 7.35 ;
      RECT  101.32 6.98 101.68 7.35 ;
      RECT  101.32 1.17 101.68 1.54 ;
      RECT  98.72 1.17 99.08 1.54 ;
      RECT  94.54 20.29 94.91 19.91 ;
      RECT  101.32 7.35 101.68 6.98 ;
      RECT  96.76 12.94 97.13 12.57 ;
      RECT  99.74 20.29 100.11 19.91 ;
      RECT  94.16 12.94 94.53 12.57 ;
      RECT  98.72 7.35 99.08 6.98 ;
      RECT  97.14 20.29 97.51 19.91 ;
      RECT  94.16 8.57 94.53 8.2 ;
      RECT  98.72 1.54 99.08 1.17 ;
      RECT  96.76 8.57 97.13 8.2 ;
      RECT  101.32 1.54 101.68 1.17 ;
      RECT  3.99 49.18 4.35 49.56 ;
      RECT  3.99 39.0 4.35 39.38 ;
      RECT  15.49 49.18 15.85 49.56 ;
      RECT  15.49 39.0 15.85 39.38 ;
      RECT  15.49 33.92 15.85 34.28 ;
      RECT  15.49 44.1 15.85 44.46 ;
      RECT  3.99 54.28 4.35 54.64 ;
      RECT  3.99 33.92 4.35 34.28 ;
      RECT  3.99 44.1 4.35 44.46 ;
      RECT  15.49 54.28 15.85 54.64 ;
      RECT  3.99 79.72 4.35 80.1 ;
      RECT  3.99 69.54 4.35 69.92 ;
      RECT  15.49 79.72 15.85 80.1 ;
      RECT  15.49 69.54 15.85 69.92 ;
      RECT  15.49 64.46 15.85 64.82 ;
      RECT  15.49 74.64 15.85 75.0 ;
      RECT  3.99 84.82 4.35 85.18 ;
      RECT  3.99 64.46 4.35 64.82 ;
      RECT  3.99 74.64 4.35 75.0 ;
      RECT  15.49 84.82 15.85 85.18 ;
      RECT  3.99 79.72 4.35 80.1 ;
      RECT  62.65 100.08 63.01 100.46 ;
      RECT  62.65 100.08 63.01 100.46 ;
      RECT  3.99 69.54 4.35 69.92 ;
      RECT  62.65 110.26 63.01 110.64 ;
      RECT  62.65 89.9 63.01 90.28 ;
      RECT  3.99 49.18 4.35 49.56 ;
      RECT  62.65 69.54 63.01 69.92 ;
      RECT  62.65 79.72 63.01 80.1 ;
      RECT  62.65 49.18 63.01 49.56 ;
      RECT  15.49 79.72 15.85 80.1 ;
      RECT  15.49 69.54 15.85 69.92 ;
      RECT  62.65 39.0 63.01 39.38 ;
      RECT  62.65 59.36 63.01 59.74 ;
      RECT  3.99 39.0 4.35 39.38 ;
      RECT  15.49 49.18 15.85 49.56 ;
      RECT  15.49 39.0 15.85 39.38 ;
      RECT  62.65 33.92 63.01 34.28 ;
      RECT  3.99 54.28 4.35 54.64 ;
      RECT  62.65 95.0 63.01 95.36 ;
      RECT  3.99 44.1 4.35 44.46 ;
      RECT  3.99 64.46 4.35 64.82 ;
      RECT  15.49 54.28 15.85 54.64 ;
      RECT  62.65 115.36 63.01 115.72 ;
      RECT  62.65 44.1 63.01 44.46 ;
      RECT  62.65 54.28 63.01 54.64 ;
      RECT  62.65 74.64 63.01 75.0 ;
      RECT  15.49 64.46 15.85 64.82 ;
      RECT  62.65 84.82 63.01 85.18 ;
      RECT  15.49 33.92 15.85 34.28 ;
      RECT  15.49 74.64 15.85 75.0 ;
      RECT  3.99 33.92 4.35 34.28 ;
      RECT  3.99 84.82 4.35 85.18 ;
      RECT  15.49 84.82 15.85 85.18 ;
      RECT  62.65 64.46 63.01 64.82 ;
      RECT  15.49 44.1 15.85 44.46 ;
      RECT  3.99 74.64 4.35 75.0 ;
      RECT  62.65 105.18 63.01 105.54 ;
      RECT  83.83 49.18 84.19 49.56 ;
      RECT  83.83 79.72 84.19 80.1 ;
      RECT  83.83 100.08 84.19 100.46 ;
      RECT  83.83 69.54 84.19 69.92 ;
      RECT  83.83 89.9 84.19 90.28 ;
      RECT  83.83 59.36 84.19 59.74 ;
      RECT  83.83 110.26 84.19 110.64 ;
      RECT  83.83 39.0 84.19 39.38 ;
      RECT  83.83 100.08 84.19 100.46 ;
      RECT  83.83 95.0 84.19 95.36 ;
      RECT  83.83 54.28 84.19 54.64 ;
      RECT  83.83 115.36 84.19 115.72 ;
      RECT  83.83 74.64 84.19 75.0 ;
      RECT  83.83 33.92 84.19 34.28 ;
      RECT  83.83 84.82 84.19 85.18 ;
      RECT  83.83 64.46 84.19 64.82 ;
      RECT  83.83 105.18 84.19 105.54 ;
      RECT  83.83 44.1 84.19 44.46 ;
      RECT  83.83 89.9 84.19 90.28 ;
      RECT  15.49 49.18 15.85 49.56 ;
      RECT  3.99 39.0 4.35 39.38 ;
      RECT  62.64 28.82 63.02 29.2 ;
      RECT  62.65 100.08 63.01 100.46 ;
      RECT  62.65 39.0 63.01 39.38 ;
      RECT  83.83 69.54 84.19 69.92 ;
      RECT  69.06 31.08 69.43 31.45 ;
      RECT  83.83 59.36 84.19 59.74 ;
      RECT  62.65 49.18 63.01 49.56 ;
      RECT  83.83 110.26 84.19 110.64 ;
      RECT  15.49 39.0 15.85 39.38 ;
      RECT  15.49 69.54 15.85 69.92 ;
      RECT  3.99 49.18 4.35 49.56 ;
      RECT  15.49 79.72 15.85 80.1 ;
      RECT  3.99 69.54 4.35 69.92 ;
      RECT  62.65 59.36 63.01 59.74 ;
      RECT  62.65 79.72 63.01 80.1 ;
      RECT  62.65 110.26 63.01 110.64 ;
      RECT  83.83 100.08 84.19 100.46 ;
      RECT  83.83 79.72 84.19 80.1 ;
      RECT  83.83 39.0 84.19 39.38 ;
      RECT  83.83 49.18 84.19 49.56 ;
      RECT  62.65 69.54 63.01 69.92 ;
      RECT  62.65 89.9 63.01 90.28 ;
      RECT  3.99 79.72 4.35 80.1 ;
      RECT  3.99 54.28 4.35 54.64 ;
      RECT  3.99 44.1 4.35 44.46 ;
      RECT  15.49 64.46 15.85 64.82 ;
      RECT  62.65 84.82 63.01 85.18 ;
      RECT  83.83 44.1 84.19 44.46 ;
      RECT  83.83 74.64 84.19 75.0 ;
      RECT  83.83 33.92 84.19 34.28 ;
      RECT  62.65 95.0 63.01 95.36 ;
      RECT  15.49 84.82 15.85 85.18 ;
      RECT  62.65 115.36 63.01 115.72 ;
      RECT  3.99 84.82 4.35 85.18 ;
      RECT  62.65 74.64 63.01 75.0 ;
      RECT  15.49 44.1 15.85 44.46 ;
      RECT  83.83 54.28 84.19 54.64 ;
      RECT  62.65 33.92 63.01 34.28 ;
      RECT  83.83 105.18 84.19 105.54 ;
      RECT  83.83 95.0 84.19 95.36 ;
      RECT  62.65 64.46 63.01 64.82 ;
      RECT  62.65 44.1 63.01 44.46 ;
      RECT  15.49 33.92 15.85 34.28 ;
      RECT  62.65 105.18 63.01 105.54 ;
      RECT  15.49 74.64 15.85 75.0 ;
      RECT  3.99 33.92 4.35 34.28 ;
      RECT  15.49 54.28 15.85 54.64 ;
      RECT  83.83 64.46 84.19 64.82 ;
      RECT  3.99 74.64 4.35 75.0 ;
      RECT  3.99 64.46 4.35 64.82 ;
      RECT  83.83 115.36 84.19 115.72 ;
      RECT  83.83 84.82 84.19 85.18 ;
      RECT  62.65 54.28 63.01 54.64 ;
      RECT  0.0 13.46 89.52 13.76 ;
      RECT  15.49 79.72 15.85 80.1 ;
      RECT  97.92 100.08 98.3 100.45 ;
      RECT  97.92 120.44 98.3 120.81 ;
      RECT  97.92 28.82 98.3 29.19 ;
      RECT  87.52 49.18 87.9 49.55 ;
      RECT  95.32 120.44 95.7 120.81 ;
      RECT  15.49 69.54 15.85 69.92 ;
      RECT  87.52 100.08 87.9 100.45 ;
      RECT  62.65 49.18 63.01 49.56 ;
      RECT  87.52 89.9 87.9 90.27 ;
      RECT  87.52 39.0 87.9 39.37 ;
      RECT  62.65 69.54 63.01 69.92 ;
      RECT  97.14 19.91 97.51 20.29 ;
      RECT  87.52 110.27 87.9 110.64 ;
      RECT  97.92 69.54 98.3 69.91 ;
      RECT  99.74 19.91 100.11 20.29 ;
      RECT  97.92 39.01 98.3 39.38 ;
      RECT  94.54 19.91 94.91 20.29 ;
      RECT  83.83 100.08 84.19 100.46 ;
      RECT  87.52 100.09 87.9 100.46 ;
      RECT  83.83 110.26 84.19 110.64 ;
      RECT  94.16 12.57 94.53 12.94 ;
      RECT  3.99 39.0 4.35 39.38 ;
      RECT  95.32 28.82 95.7 29.19 ;
      RECT  101.32 6.98 101.68 7.35 ;
      RECT  97.92 59.37 98.3 59.74 ;
      RECT  97.92 110.26 98.3 110.63 ;
      RECT  97.92 69.55 98.3 69.92 ;
      RECT  87.52 89.91 87.9 90.28 ;
      RECT  83.83 39.0 84.19 39.38 ;
      RECT  69.06 31.08 69.43 31.45 ;
      RECT  3.99 49.18 4.35 49.56 ;
      RECT  62.65 79.72 63.01 80.1 ;
      RECT  87.52 110.26 87.9 110.63 ;
      RECT  62.65 39.0 63.01 39.38 ;
      RECT  83.83 89.9 84.19 90.28 ;
      RECT  83.83 49.18 84.19 49.56 ;
      RECT  87.52 49.19 87.9 49.56 ;
      RECT  15.49 49.18 15.85 49.56 ;
      RECT  62.64 28.82 63.02 29.2 ;
      RECT  83.83 79.72 84.19 80.1 ;
      RECT  15.49 39.0 15.85 39.38 ;
      RECT  87.52 28.82 87.9 29.19 ;
      RECT  90.13 28.82 90.49 29.19 ;
      RECT  97.92 100.09 98.3 100.46 ;
      RECT  87.52 69.54 87.9 69.91 ;
      RECT  92.72 28.82 93.1 29.19 ;
      RECT  97.92 79.73 98.3 80.1 ;
      RECT  97.92 89.9 98.3 90.27 ;
      RECT  3.99 79.72 4.35 80.1 ;
      RECT  62.65 59.36 63.01 59.74 ;
      RECT  97.92 110.27 98.3 110.64 ;
      RECT  83.83 69.54 84.19 69.92 ;
      RECT  97.92 28.83 98.3 29.2 ;
      RECT  92.72 120.44 93.1 120.81 ;
      RECT  97.92 39.0 98.3 39.37 ;
      RECT  87.52 79.72 87.9 80.09 ;
      RECT  62.65 100.08 63.01 100.46 ;
      RECT  3.99 69.54 4.35 69.92 ;
      RECT  96.76 12.57 97.13 12.94 ;
      RECT  87.52 120.44 87.9 120.81 ;
      RECT  87.52 79.73 87.9 80.1 ;
      RECT  83.83 59.36 84.19 59.74 ;
      RECT  97.92 49.19 98.3 49.56 ;
      RECT  62.65 89.9 63.01 90.28 ;
      RECT  87.52 59.36 87.9 59.73 ;
      RECT  87.52 39.01 87.9 39.38 ;
      RECT  87.52 69.55 87.9 69.92 ;
      RECT  98.72 6.98 99.08 7.35 ;
      RECT  87.52 59.37 87.9 59.74 ;
      RECT  97.92 79.72 98.3 80.09 ;
      RECT  97.92 59.36 98.3 59.73 ;
      RECT  97.92 89.91 98.3 90.28 ;
      RECT  90.13 120.44 90.49 120.81 ;
      RECT  62.65 110.26 63.01 110.64 ;
      RECT  97.92 49.18 98.3 49.55 ;
      RECT  87.52 28.83 87.9 29.2 ;
      RECT  101.32 1.17 101.68 1.54 ;
      RECT  83.83 44.1 84.19 44.46 ;
      RECT  62.65 64.46 63.01 64.82 ;
      RECT  97.92 44.09 98.3 44.46 ;
      RECT  99.92 24.88 100.28 25.26 ;
      RECT  83.83 115.36 84.19 115.72 ;
      RECT  3.99 84.82 4.35 85.18 ;
      RECT  15.49 33.92 15.85 34.28 ;
      RECT  3.99 33.92 4.35 34.28 ;
      RECT  85.54 24.88 85.9 25.26 ;
      RECT  15.49 84.82 15.85 85.18 ;
      RECT  62.65 84.82 63.01 85.18 ;
      RECT  95.32 23.74 95.7 24.11 ;
      RECT  97.92 44.1 98.3 44.47 ;
      RECT  87.52 64.46 87.9 64.83 ;
      RECT  90.13 115.36 90.49 115.73 ;
      RECT  15.49 74.64 15.85 75.0 ;
      RECT  87.52 74.64 87.9 75.01 ;
      RECT  87.52 105.17 87.9 105.54 ;
      RECT  97.92 115.35 98.3 115.72 ;
      RECT  87.52 54.27 87.9 54.64 ;
      RECT  85.54 116.5 85.9 116.88 ;
      RECT  87.52 33.92 87.9 34.29 ;
      RECT  97.92 74.63 98.3 75.0 ;
      RECT  62.65 33.92 63.01 34.28 ;
      RECT  83.83 84.82 84.19 85.18 ;
      RECT  62.65 74.64 63.01 75.0 ;
      RECT  99.92 116.5 100.28 116.88 ;
      RECT  97.92 54.28 98.3 54.65 ;
      RECT  87.52 105.18 87.9 105.55 ;
      RECT  62.65 105.18 63.01 105.54 ;
      RECT  87.52 44.1 87.9 44.47 ;
      RECT  90.13 23.74 90.49 24.11 ;
      RECT  97.92 105.17 98.3 105.54 ;
      RECT  97.92 95.0 98.3 95.37 ;
      RECT  97.92 84.81 98.3 85.18 ;
      RECT  87.52 115.36 87.9 115.73 ;
      RECT  97.92 94.99 98.3 95.36 ;
      RECT  97.92 23.74 98.3 24.11 ;
      RECT  3.99 44.1 4.35 44.46 ;
      RECT  97.92 64.46 98.3 64.83 ;
      RECT  97.92 33.92 98.3 34.29 ;
      RECT  83.83 33.92 84.19 34.28 ;
      RECT  87.52 94.99 87.9 95.36 ;
      RECT  97.92 64.45 98.3 64.82 ;
      RECT  62.65 54.28 63.01 54.64 ;
      RECT  96.76 8.2 97.13 8.57 ;
      RECT  94.16 8.2 94.53 8.57 ;
      RECT  98.72 1.17 99.08 1.54 ;
      RECT  87.52 74.63 87.9 75.0 ;
      RECT  3.99 64.46 4.35 64.82 ;
      RECT  87.52 33.91 87.9 34.28 ;
      RECT  83.83 74.64 84.19 75.0 ;
      RECT  97.92 74.64 98.3 75.01 ;
      RECT  15.49 54.28 15.85 54.64 ;
      RECT  87.52 54.28 87.9 54.65 ;
      RECT  83.83 54.28 84.19 54.64 ;
      RECT  87.52 95.0 87.9 95.37 ;
      RECT  15.49 44.1 15.85 44.46 ;
      RECT  87.52 115.35 87.9 115.72 ;
      RECT  3.99 74.64 4.35 75.0 ;
      RECT  83.83 64.46 84.19 64.82 ;
      RECT  62.65 95.0 63.01 95.36 ;
      RECT  3.99 54.28 4.35 54.64 ;
      RECT  97.92 84.82 98.3 85.19 ;
      RECT  83.83 95.0 84.19 95.36 ;
      RECT  92.72 23.74 93.1 24.11 ;
      RECT  97.92 105.18 98.3 105.55 ;
      RECT  87.52 64.45 87.9 64.82 ;
      RECT  87.52 84.81 87.9 85.18 ;
      RECT  95.32 115.36 95.7 115.73 ;
      RECT  97.92 115.36 98.3 115.73 ;
      RECT  97.92 33.91 98.3 34.28 ;
      RECT  87.52 23.74 87.9 24.11 ;
      RECT  97.92 54.27 98.3 54.64 ;
      RECT  87.52 44.09 87.9 44.46 ;
      RECT  62.65 115.36 63.01 115.72 ;
      RECT  62.65 44.1 63.01 44.46 ;
      RECT  15.49 64.46 15.85 64.82 ;
      RECT  92.72 115.36 93.1 115.73 ;
      RECT  83.83 105.18 84.19 105.54 ;
      RECT  87.52 84.82 87.9 85.19 ;
      RECT  -103.49 -5.61 -103.13 -5.24 ;
      RECT  -103.49 -5.6 -103.13 -5.23 ;
      RECT  -103.55 -9.69 -103.19 -9.32 ;
      RECT  -103.55 -1.52 -103.19 -1.15 ;
      RECT  -93.23 43.06 -93.59 43.42 ;
      RECT  -76.35 55.94 -76.71 56.3 ;
      RECT  -93.23 68.82 -93.59 69.18 ;
      RECT  -76.35 81.7 -76.71 82.06 ;
      RECT  -93.23 55.94 -93.59 56.3 ;
      RECT  -76.35 43.06 -76.71 43.42 ;
      RECT  -76.35 30.18 -76.71 30.54 ;
      RECT  -93.23 81.7 -93.59 82.06 ;
      RECT  -93.23 30.18 -93.59 30.54 ;
      RECT  -76.35 68.82 -76.71 69.18 ;
      RECT  -93.23 36.62 -93.59 36.98 ;
      RECT  -76.35 62.38 -76.71 62.74 ;
      RECT  -76.35 36.62 -76.71 36.98 ;
      RECT  -76.35 75.26 -76.71 75.62 ;
      RECT  -93.23 75.26 -93.59 75.62 ;
      RECT  -76.35 23.74 -76.71 24.1 ;
      RECT  -93.23 49.5 -93.59 49.86 ;
      RECT  -76.35 49.5 -76.71 49.86 ;
      RECT  -93.23 23.74 -93.59 24.1 ;
      RECT  -93.23 62.38 -93.59 62.74 ;
      RECT  -93.59 55.94 -93.23 56.3 ;
      RECT  -76.71 30.18 -76.35 30.54 ;
      RECT  -103.49 -5.6 -103.13 -5.23 ;
      RECT  -76.71 68.82 -76.35 69.18 ;
      RECT  -93.59 30.18 -93.23 30.54 ;
      RECT  -76.71 43.06 -76.35 43.42 ;
      RECT  -93.59 43.06 -93.23 43.42 ;
      RECT  -103.49 -5.61 -103.13 -5.24 ;
      RECT  -93.59 68.82 -93.23 69.18 ;
      RECT  -76.71 81.7 -76.35 82.06 ;
      RECT  -93.59 81.7 -93.23 82.06 ;
      RECT  -76.71 55.94 -76.35 56.3 ;
      RECT  -93.59 49.5 -93.23 49.86 ;
      RECT  -76.71 62.38 -76.35 62.74 ;
      RECT  -76.71 49.5 -76.35 49.86 ;
      RECT  -76.71 36.62 -76.35 36.98 ;
      RECT  -76.71 75.26 -76.35 75.62 ;
      RECT  -93.59 36.62 -93.23 36.98 ;
      RECT  -103.55 -9.69 -103.19 -9.32 ;
      RECT  -76.71 23.74 -76.35 24.1 ;
      RECT  -93.59 62.38 -93.23 62.74 ;
      RECT  -93.59 23.74 -93.23 24.1 ;
      RECT  -93.59 75.26 -93.23 75.62 ;
      RECT  -103.55 -1.52 -103.19 -1.15 ;
      RECT  -12.67 84.31 -1.02 84.61 ;
      RECT  -7.53 86.67 -7.16 87.04 ;
      RECT  -7.53 94.79 -7.16 95.16 ;
      RECT  -7.53 94.8 -7.16 95.17 ;
      RECT  -7.53 86.68 -7.16 87.05 ;
      RECT  -7.65 98.88 -7.28 99.25 ;
      RECT  -7.65 90.76 -7.28 91.13 ;
      RECT  -7.65 82.59 -7.28 82.96 ;
      RECT  -7.65 90.71 -7.28 91.08 ;
      RECT  10.63 -7.97 33.93 -7.67 ;
      RECT  27.42 -5.6 27.79 -5.23 ;
      RECT  15.77 -5.6 16.14 -5.23 ;
      RECT  15.65 -9.69 16.02 -9.32 ;
      RECT  27.3 -9.69 27.67 -9.32 ;
   LAYER  m4 ;
   END
   END    sram_2_16_sky130A
END    LIBRARY
