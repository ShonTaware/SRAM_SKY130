magic
tech sky130A
timestamp 1613393220
<< fence >>
rect 155 -252 913 425
<< nwell >>
rect 170 -22 327 198
rect 455 -44 735 210
rect 455 -45 657 -44
<< nmos >>
rect 259 317 274 359
rect 520 317 535 359
rect 664 317 679 359
rect 805 317 820 359
rect 259 -179 274 -137
rect 512 -180 527 -138
rect 664 -180 679 -138
rect 803 -180 818 -138
<< pmos >>
rect 259 138 274 180
rect 259 -4 274 38
rect 520 148 535 190
rect 664 148 679 190
rect 512 -25 527 17
rect 664 -25 679 17
<< ndiff >>
rect 220 350 259 359
rect 220 333 226 350
rect 243 333 259 350
rect 220 317 259 333
rect 274 348 314 359
rect 274 331 288 348
rect 305 331 314 348
rect 274 317 314 331
rect 480 348 520 359
rect 480 329 484 348
rect 503 329 520 348
rect 480 317 520 329
rect 535 348 576 359
rect 535 329 551 348
rect 570 329 576 348
rect 535 317 576 329
rect 617 346 664 359
rect 617 327 623 346
rect 642 327 664 346
rect 617 317 664 327
rect 679 349 735 359
rect 679 330 709 349
rect 728 330 735 349
rect 679 317 735 330
rect 764 347 805 359
rect 764 328 769 347
rect 788 328 805 347
rect 764 317 805 328
rect 820 345 861 359
rect 820 326 836 345
rect 855 326 861 345
rect 820 317 861 326
rect 220 -153 259 -137
rect 220 -170 226 -153
rect 243 -170 259 -153
rect 220 -179 259 -170
rect 274 -151 314 -137
rect 274 -168 288 -151
rect 305 -168 314 -151
rect 274 -179 314 -168
rect 474 -147 512 -138
rect 474 -169 479 -147
rect 497 -169 512 -147
rect 474 -180 512 -169
rect 527 -148 565 -138
rect 527 -170 543 -148
rect 561 -170 565 -148
rect 527 -180 565 -170
rect 620 -148 664 -138
rect 620 -170 626 -148
rect 644 -170 664 -148
rect 620 -180 664 -170
rect 679 -147 723 -138
rect 679 -169 695 -147
rect 713 -169 723 -147
rect 679 -180 723 -169
rect 761 -149 803 -138
rect 761 -169 767 -149
rect 784 -169 803 -149
rect 761 -180 803 -169
rect 818 -146 863 -138
rect 818 -168 841 -146
rect 859 -168 863 -146
rect 818 -180 863 -168
<< pdiff >>
rect 224 171 259 180
rect 224 148 229 171
rect 246 148 259 171
rect 224 138 259 148
rect 274 171 309 180
rect 274 148 288 171
rect 305 148 309 171
rect 274 138 309 148
rect 224 28 259 38
rect 224 5 229 28
rect 246 5 259 28
rect 224 -4 259 5
rect 274 28 309 38
rect 274 5 288 28
rect 305 5 309 28
rect 274 -4 309 5
rect 485 182 520 190
rect 485 159 489 182
rect 506 159 520 182
rect 485 148 520 159
rect 535 179 570 190
rect 535 156 548 179
rect 565 156 570 179
rect 535 148 570 156
rect 627 182 664 190
rect 627 159 634 182
rect 651 159 664 182
rect 627 148 664 159
rect 679 182 716 190
rect 679 159 694 182
rect 711 159 716 182
rect 679 148 716 159
rect 479 6 512 17
rect 479 -17 483 6
rect 500 -17 512 6
rect 479 -25 512 -17
rect 527 9 560 17
rect 527 -14 536 9
rect 553 -14 560 9
rect 527 -25 560 -14
rect 627 6 664 17
rect 627 -17 633 6
rect 650 -17 664 6
rect 627 -25 664 -17
rect 679 6 716 17
rect 679 -17 694 6
rect 711 -17 716 6
rect 679 -25 716 -17
<< ndiffc >>
rect 226 333 243 350
rect 288 331 305 348
rect 484 329 503 348
rect 551 329 570 348
rect 623 327 642 346
rect 709 330 728 349
rect 769 328 788 347
rect 836 326 855 345
rect 226 -170 243 -153
rect 288 -168 305 -151
rect 479 -169 497 -147
rect 543 -170 561 -148
rect 626 -170 644 -148
rect 695 -169 713 -147
rect 767 -169 784 -149
rect 841 -168 859 -146
<< pdiffc >>
rect 229 148 246 171
rect 288 148 305 171
rect 229 5 246 28
rect 288 5 305 28
rect 489 159 506 182
rect 548 156 565 179
rect 634 159 651 182
rect 694 159 711 182
rect 483 -17 500 6
rect 536 -14 553 9
rect 633 -17 650 6
rect 694 -17 711 6
<< psubdiff >>
rect 202 396 256 422
rect 287 396 517 422
rect 548 396 653 422
rect 684 396 753 422
rect 784 396 811 422
rect 466 395 486 396
rect 202 -242 256 -216
rect 287 -242 341 -216
rect 547 -217 613 -208
rect 709 -217 728 -210
rect 457 -243 511 -217
rect 542 -243 653 -217
rect 684 -243 733 -217
rect 764 -243 808 -217
rect 547 -244 613 -243
<< nsubdiff >>
rect 222 84 241 85
rect 202 65 245 84
rect 268 65 309 84
rect 473 66 487 85
rect 504 66 531 85
<< psubdiffcont >>
rect 256 396 287 422
rect 517 396 548 422
rect 653 396 684 422
rect 753 396 784 422
rect 256 -242 287 -216
rect 511 -243 542 -217
rect 653 -243 684 -217
rect 733 -243 764 -217
<< nsubdiffcont >>
rect 245 65 268 84
rect 487 66 504 85
<< poly >>
rect 259 359 274 372
rect 520 359 535 372
rect 664 359 679 372
rect 805 359 820 372
rect 259 232 274 317
rect 432 286 470 296
rect 520 286 535 317
rect 432 285 535 286
rect 432 266 442 285
rect 460 271 535 285
rect 460 266 470 271
rect 432 258 470 266
rect 259 217 375 232
rect 259 180 274 217
rect 259 125 274 138
rect 259 38 274 51
rect 259 -51 274 -4
rect 176 -61 274 -51
rect 176 -83 183 -61
rect 203 -83 274 -61
rect 360 -68 375 217
rect 520 190 535 271
rect 664 190 679 317
rect 805 292 820 317
rect 796 284 834 292
rect 796 265 806 284
rect 824 265 834 284
rect 796 254 834 265
rect 520 135 535 148
rect 664 97 679 148
rect 761 100 797 112
rect 761 97 768 100
rect 664 82 768 97
rect 512 17 527 30
rect 664 17 679 82
rect 761 77 768 82
rect 788 77 797 100
rect 761 65 797 77
rect 176 -93 274 -83
rect 259 -137 274 -93
rect 352 -78 390 -68
rect 352 -97 360 -78
rect 378 -81 390 -78
rect 512 -81 527 -25
rect 378 -96 527 -81
rect 378 -97 390 -96
rect 352 -106 390 -97
rect 512 -138 527 -96
rect 664 -138 679 -25
rect 787 -70 825 -62
rect 787 -89 797 -70
rect 815 -89 825 -70
rect 787 -100 825 -89
rect 803 -138 818 -100
rect 259 -192 274 -179
rect 512 -193 527 -180
rect 664 -193 679 -180
rect 803 -193 818 -180
<< polycont >>
rect 442 266 460 285
rect 183 -83 203 -61
rect 806 265 824 284
rect 768 77 788 100
rect 360 -97 378 -78
rect 797 -89 815 -70
<< locali >>
rect 195 422 812 423
rect 195 396 256 422
rect 287 415 517 422
rect 287 396 466 415
rect 486 396 517 415
rect 548 396 653 422
rect 684 416 753 422
rect 684 397 717 416
rect 737 397 753 416
rect 684 396 753 397
rect 784 416 812 422
rect 784 397 790 416
rect 810 397 812 416
rect 784 396 812 397
rect 195 394 812 396
rect 227 359 244 394
rect 486 359 504 394
rect 623 359 640 394
rect 769 359 786 394
rect 220 350 252 359
rect 220 333 226 350
rect 243 333 252 350
rect 220 323 252 333
rect 282 348 314 359
rect 282 331 288 348
rect 305 331 314 348
rect 282 323 314 331
rect 480 348 509 359
rect 480 329 484 348
rect 503 329 509 348
rect 289 286 306 323
rect 480 317 509 329
rect 547 348 576 359
rect 547 329 551 348
rect 570 329 576 348
rect 547 317 576 329
rect 617 346 646 359
rect 617 327 623 346
rect 642 327 646 346
rect 617 317 646 327
rect 702 349 731 359
rect 702 330 709 349
rect 728 330 731 349
rect 702 317 731 330
rect 764 347 793 359
rect 764 328 769 347
rect 788 328 793 347
rect 764 317 793 328
rect 832 345 861 359
rect 832 326 836 345
rect 855 343 861 345
rect 855 326 887 343
rect 904 326 907 343
rect 832 317 861 326
rect 432 286 470 296
rect 289 285 470 286
rect 289 269 442 285
rect 289 179 306 269
rect 432 266 442 269
rect 460 266 470 285
rect 432 258 470 266
rect 553 282 570 317
rect 707 282 724 317
rect 796 284 834 292
rect 796 282 806 284
rect 553 265 806 282
rect 824 265 834 284
rect 695 190 712 265
rect 796 254 834 265
rect 485 182 512 190
rect 224 171 251 179
rect 224 148 229 171
rect 246 148 251 171
rect 224 138 251 148
rect 282 171 309 179
rect 282 148 288 171
rect 305 148 309 171
rect 485 159 489 182
rect 506 159 512 182
rect 485 149 512 159
rect 543 179 570 190
rect 543 156 548 179
rect 565 178 570 179
rect 627 182 654 190
rect 627 178 634 182
rect 565 161 634 178
rect 565 156 570 161
rect 282 138 309 148
rect 228 87 245 138
rect 492 88 509 149
rect 543 148 570 156
rect 627 159 634 161
rect 651 159 654 182
rect 627 148 654 159
rect 689 182 716 190
rect 689 159 694 182
rect 711 159 716 182
rect 689 149 716 159
rect 761 100 797 112
rect 197 61 200 87
rect 221 84 291 87
rect 221 65 245 84
rect 268 65 291 84
rect 221 61 291 65
rect 312 61 316 87
rect 473 85 548 88
rect 473 66 487 85
rect 504 82 548 85
rect 504 66 524 82
rect 473 65 524 66
rect 541 65 548 82
rect 761 77 768 100
rect 788 98 797 100
rect 788 81 814 98
rect 788 77 797 81
rect 761 65 797 77
rect 473 62 548 65
rect 228 38 245 61
rect 224 28 251 38
rect 224 5 229 28
rect 246 5 251 28
rect 224 -3 251 5
rect 282 28 309 38
rect 282 5 288 28
rect 305 5 309 28
rect 483 16 500 62
rect 282 -3 309 5
rect 479 6 506 16
rect 176 -61 211 -51
rect 176 -66 183 -61
rect 155 -83 183 -66
rect 203 -83 211 -61
rect 176 -93 211 -83
rect 289 -79 306 -3
rect 479 -17 483 6
rect 500 -17 506 6
rect 479 -25 506 -17
rect 533 9 560 17
rect 533 -14 536 9
rect 553 6 560 9
rect 627 6 654 17
rect 553 -11 633 6
rect 553 -14 560 -11
rect 533 -25 560 -14
rect 627 -17 633 -11
rect 650 -17 654 6
rect 627 -25 654 -17
rect 689 6 716 16
rect 689 -17 694 6
rect 711 -17 716 6
rect 689 -25 716 -17
rect 352 -78 390 -68
rect 695 -73 712 -25
rect 787 -70 825 -62
rect 787 -73 797 -70
rect 352 -79 360 -78
rect 289 -96 360 -79
rect 289 -143 306 -96
rect 352 -97 360 -96
rect 378 -97 390 -78
rect 352 -106 390 -97
rect 543 -89 797 -73
rect 815 -89 825 -70
rect 543 -90 825 -89
rect 543 -138 560 -90
rect 695 -138 712 -90
rect 787 -100 825 -90
rect 220 -153 252 -143
rect 220 -170 226 -153
rect 243 -170 252 -153
rect 220 -179 252 -170
rect 282 -151 314 -143
rect 282 -168 288 -151
rect 305 -168 314 -151
rect 282 -179 314 -168
rect 474 -147 503 -138
rect 474 -169 479 -147
rect 497 -169 503 -147
rect 227 -208 244 -179
rect 474 -180 503 -169
rect 536 -148 565 -138
rect 536 -170 543 -148
rect 561 -170 565 -148
rect 536 -180 565 -170
rect 620 -148 649 -138
rect 620 -170 626 -148
rect 644 -170 649 -148
rect 620 -180 649 -170
rect 689 -147 718 -138
rect 689 -169 695 -147
rect 713 -169 718 -147
rect 689 -180 718 -169
rect 761 -149 792 -138
rect 761 -169 767 -149
rect 784 -169 792 -149
rect 761 -180 792 -169
rect 832 -146 863 -138
rect 832 -168 841 -146
rect 859 -152 863 -146
rect 859 -168 891 -152
rect 832 -169 891 -168
rect 832 -180 863 -169
rect 195 -209 424 -208
rect 480 -209 498 -180
rect 624 -208 641 -180
rect 543 -209 650 -208
rect 696 -209 713 -208
rect 770 -209 787 -180
rect 195 -216 826 -209
rect 195 -233 224 -216
rect 241 -233 256 -216
rect 195 -242 256 -233
rect 287 -217 826 -216
rect 287 -218 511 -217
rect 287 -235 460 -218
rect 477 -235 511 -218
rect 287 -242 511 -235
rect 195 -243 511 -242
rect 542 -220 653 -217
rect 542 -237 588 -220
rect 605 -237 653 -220
rect 542 -243 653 -237
rect 684 -243 733 -217
rect 764 -243 777 -217
rect 808 -243 826 -217
rect 448 -244 826 -243
<< viali >>
rect 466 396 486 415
rect 717 397 737 416
rect 790 397 810 416
rect 887 326 904 343
rect 200 61 221 87
rect 291 61 312 87
rect 524 65 541 82
rect 891 -169 908 -152
rect 224 -233 241 -216
rect 460 -235 477 -218
rect 588 -237 605 -220
rect 777 -243 808 -217
<< metal1 >>
rect 193 416 814 425
rect 193 415 717 416
rect 193 396 466 415
rect 486 397 717 415
rect 737 397 790 416
rect 810 397 814 416
rect 486 396 814 397
rect 193 387 814 396
rect 861 343 910 351
rect 861 326 887 343
rect 904 326 910 343
rect 861 320 910 326
rect 188 87 320 95
rect 188 61 200 87
rect 221 61 291 87
rect 312 61 320 87
rect 188 54 320 61
rect 455 82 548 96
rect 455 65 524 82
rect 541 65 548 82
rect 455 55 548 65
rect 863 -152 913 -146
rect 863 -169 891 -152
rect 908 -169 913 -152
rect 863 -174 913 -169
rect 899 -175 913 -174
rect 185 -208 244 -207
rect 185 -216 826 -208
rect 185 -233 224 -216
rect 241 -217 826 -216
rect 241 -218 777 -217
rect 241 -233 460 -218
rect 185 -235 460 -233
rect 477 -220 777 -218
rect 477 -235 588 -220
rect 185 -237 588 -235
rect 605 -237 777 -220
rect 185 -243 777 -237
rect 808 -243 826 -217
rect 185 -252 826 -243
<< labels >>
flabel locali 308 -96 331 -80 0 FreeSans 80 0 0 0 dinb
flabel metal1 224 63 243 80 0 FreeSans 72 270 0 0 vdd
flabel metal1 507 65 520 82 0 FreeSans 72 270 0 0 vdd
flabel metal1 559 395 613 422 0 FreeSans 152 0 0 0 gnd
flabel metal1 294 -242 341 -216 0 FreeSans 152 0 0 0 gnd
flabel locali 291 270 346 285 0 FreeSans 152 0 0 0 dinbb
flabel locali 156 -82 175 -67 0 FreeSans 120 0 0 0 din
flabel locali 704 -89 745 -73 0 FreeSans 144 0 0 0 out1
flabel locali 707 266 739 282 0 FreeSans 144 0 0 0 out2
flabel metal1 863 327 886 343 0 FreeSans 120 0 0 0 bl
flabel metal1 866 -167 888 -153 0 FreeSans 96 0 0 0 blbar
flabel locali 575 -10 605 5 0 FreeSans 120 0 0 0 4
flabel locali 579 162 607 177 0 FreeSans 120 0 0 0 5
flabel locali 799 83 812 95 0 FreeSans 88 0 0 0 wen
<< end >>
