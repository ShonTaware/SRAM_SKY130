magic
tech sky130A
timestamp 1615133568
<< error_p >>
rect 297 -40 298 -23
rect 316 -40 317 -23
rect 433 -40 434 -23
rect 452 -40 453 -23
<< nwell >>
rect -3 226 577 452
rect 300 225 577 226
<< nmos >>
rect 60 20 75 62
rect 230 20 245 62
rect 364 20 379 120
rect 502 20 517 62
<< pmos >>
rect 60 246 75 301
rect 230 246 245 346
rect 502 246 517 301
<< ndiff >>
rect 319 110 364 120
rect 319 93 332 110
rect 349 93 364 110
rect 15 50 60 62
rect 15 33 28 50
rect 45 33 60 50
rect 15 20 60 33
rect 75 50 115 62
rect 75 33 88 50
rect 105 33 115 50
rect 75 20 115 33
rect 185 50 230 62
rect 185 33 198 50
rect 215 33 230 50
rect 185 20 230 33
rect 245 50 285 62
rect 245 33 258 50
rect 275 33 285 50
rect 245 20 285 33
rect 319 50 364 93
rect 319 33 332 50
rect 349 33 364 50
rect 319 20 364 33
rect 379 110 419 120
rect 379 93 392 110
rect 409 93 419 110
rect 379 50 419 93
rect 379 33 392 50
rect 409 33 419 50
rect 379 20 419 33
rect 457 50 502 62
rect 457 33 470 50
rect 487 33 502 50
rect 457 20 502 33
rect 517 50 557 62
rect 517 33 530 50
rect 547 33 557 50
rect 517 20 557 33
<< pdiff >>
rect 185 335 230 346
rect 185 318 198 335
rect 215 318 230 335
rect 15 282 60 301
rect 15 265 28 282
rect 45 265 60 282
rect 15 246 60 265
rect 75 282 115 301
rect 75 265 88 282
rect 105 265 115 282
rect 75 246 115 265
rect 185 282 230 318
rect 185 265 198 282
rect 215 265 230 282
rect 185 246 230 265
rect 245 335 285 346
rect 245 318 258 335
rect 275 318 285 335
rect 245 282 285 318
rect 245 265 258 282
rect 275 265 285 282
rect 245 246 285 265
rect 457 282 502 301
rect 457 265 470 282
rect 487 265 502 282
rect 457 246 502 265
rect 517 282 557 301
rect 517 265 530 282
rect 547 265 557 282
rect 517 246 557 265
<< ndiffc >>
rect 332 93 349 110
rect 28 33 45 50
rect 88 33 105 50
rect 198 33 215 50
rect 258 33 275 50
rect 332 33 349 50
rect 392 93 409 110
rect 392 33 409 50
rect 470 33 487 50
rect 530 33 547 50
<< pdiffc >>
rect 198 318 215 335
rect 28 265 45 282
rect 88 265 105 282
rect 198 265 215 282
rect 258 318 275 335
rect 258 265 275 282
rect 470 265 487 282
rect 530 265 547 282
<< psubdiff >>
rect 48 -23 89 -11
rect 48 -40 60 -23
rect 77 -40 89 -23
rect 48 -52 89 -40
rect 218 -23 259 -11
rect 218 -40 230 -23
rect 247 -40 259 -23
rect 218 -52 259 -40
rect 354 -23 395 -11
rect 354 -40 366 -23
rect 383 -40 395 -23
rect 354 -52 395 -40
rect 490 -23 531 -11
rect 490 -40 502 -23
rect 519 -40 531 -23
rect 490 -52 531 -40
<< nsubdiff >>
rect 37 414 90 432
rect 37 397 55 414
rect 72 397 90 414
rect 37 379 90 397
rect 207 414 260 432
rect 207 397 225 414
rect 242 397 260 414
rect 207 379 260 397
rect 343 414 396 432
rect 343 397 361 414
rect 378 397 396 414
rect 343 379 396 397
rect 479 414 532 432
rect 479 397 497 414
rect 514 397 532 414
rect 479 379 532 397
<< psubdiffcont >>
rect 60 -40 77 -23
rect 230 -40 247 -23
rect 366 -40 383 -23
rect 502 -40 519 -23
<< nsubdiffcont >>
rect 55 397 72 414
rect 225 397 242 414
rect 361 397 378 414
rect 497 397 514 414
<< poly >>
rect 230 346 245 363
rect 60 301 75 318
rect 502 301 517 318
rect 60 201 75 246
rect 97 203 130 211
rect 97 201 105 203
rect 60 186 105 201
rect 122 201 130 203
rect 230 201 245 246
rect 502 215 517 246
rect 122 186 245 201
rect 439 207 517 215
rect 439 190 447 207
rect 464 200 517 207
rect 464 190 472 200
rect 97 178 130 186
rect 439 182 472 190
rect 364 130 473 145
rect 364 120 379 130
rect -29 105 4 113
rect -29 88 -21 105
rect -4 95 4 105
rect 135 105 168 113
rect -4 88 75 95
rect -29 80 75 88
rect 135 88 143 105
rect 160 95 168 105
rect 160 88 245 95
rect 135 80 245 88
rect 60 62 75 80
rect 230 62 245 80
rect 458 108 473 130
rect 445 100 478 108
rect 445 83 453 100
rect 470 83 478 100
rect 445 75 478 83
rect 502 62 517 200
rect 60 5 75 20
rect 230 5 245 20
rect 364 5 379 20
rect 502 5 517 20
<< polycont >>
rect 105 186 122 203
rect 447 190 464 207
rect -21 88 -4 105
rect 143 88 160 105
rect 453 83 470 100
<< locali >>
rect -2 414 577 422
rect -2 397 5 414
rect 22 397 55 414
rect 72 397 100 414
rect 117 397 175 414
rect 192 397 225 414
rect 242 397 270 414
rect 287 397 311 414
rect 328 397 361 414
rect 378 397 406 414
rect 423 397 447 414
rect 464 397 497 414
rect 514 397 542 414
rect 559 397 577 414
rect -2 389 577 397
rect 25 290 45 389
rect 195 343 215 389
rect 190 335 223 343
rect 190 318 198 335
rect 215 318 223 335
rect 20 282 53 290
rect 20 265 28 282
rect 45 265 53 282
rect 20 257 53 265
rect 80 282 115 290
rect 80 265 88 282
rect 105 265 115 282
rect 80 257 115 265
rect 190 282 223 318
rect 190 265 198 282
rect 215 265 223 282
rect 190 257 223 265
rect 250 335 283 343
rect 250 318 258 335
rect 275 318 283 335
rect 250 282 283 318
rect 467 290 487 389
rect 250 265 258 282
rect 275 265 283 282
rect 250 257 283 265
rect 462 282 495 290
rect 462 265 470 282
rect 487 265 495 282
rect 462 257 495 265
rect 522 282 555 290
rect 522 265 530 282
rect 547 265 555 282
rect 522 257 555 265
rect 97 211 115 257
rect 259 215 279 257
rect 97 203 130 211
rect 97 186 105 203
rect 122 186 130 203
rect 97 178 130 186
rect 259 207 472 215
rect 259 195 447 207
rect 17 168 46 174
rect 17 151 23 168
rect 40 151 46 168
rect 17 145 46 151
rect -29 105 4 113
rect -29 88 -21 105
rect -4 88 4 105
rect -29 80 4 88
rect 26 58 46 145
rect 97 58 115 178
rect 189 168 218 174
rect 189 151 195 168
rect 212 151 218 168
rect 189 145 218 151
rect 135 105 168 113
rect 135 88 143 105
rect 160 88 168 105
rect 135 80 168 88
rect 194 58 214 145
rect 259 58 279 195
rect 439 190 447 195
rect 464 190 472 207
rect 439 182 472 190
rect 315 168 344 174
rect 315 151 321 168
rect 338 151 344 168
rect 315 145 344 151
rect 324 118 344 145
rect 529 172 549 257
rect 529 166 558 172
rect 529 149 535 166
rect 552 149 558 166
rect 529 142 558 149
rect 324 110 357 118
rect 324 93 332 110
rect 349 93 357 110
rect 26 55 53 58
rect 20 50 53 55
rect 20 33 28 50
rect 45 33 53 50
rect 20 25 53 33
rect 80 50 115 58
rect 80 33 88 50
rect 105 33 115 50
rect 80 25 115 33
rect 190 50 223 58
rect 190 33 198 50
rect 215 33 223 50
rect 190 25 223 33
rect 250 50 283 58
rect 250 33 258 50
rect 275 33 283 50
rect 250 25 283 33
rect 324 50 357 93
rect 324 33 332 50
rect 349 33 357 50
rect 324 25 357 33
rect 384 110 417 118
rect 384 93 392 110
rect 409 93 417 110
rect 384 50 417 93
rect 445 100 478 108
rect 445 83 453 100
rect 470 83 478 100
rect 445 75 478 83
rect 529 58 549 142
rect 384 33 392 50
rect 409 33 417 50
rect 384 25 417 33
rect 462 50 495 58
rect 462 33 470 50
rect 487 33 495 50
rect 462 25 495 33
rect 522 50 555 58
rect 522 33 530 50
rect 547 33 555 50
rect 522 25 555 33
rect 394 -15 414 25
rect 464 -15 484 25
rect -3 -23 577 -15
rect -3 -40 10 -23
rect 27 -40 60 -23
rect 77 -40 110 -23
rect 127 -40 184 -23
rect 201 -40 230 -23
rect 247 -40 281 -23
rect 298 -40 316 -23
rect 333 -40 366 -23
rect 383 -40 417 -23
rect 434 -40 452 -23
rect 469 -40 502 -23
rect 519 -40 553 -23
rect 570 -40 577 -23
rect -3 -48 577 -40
<< viali >>
rect 5 397 22 414
rect 100 397 117 414
rect 175 397 192 414
rect 270 397 287 414
rect 311 397 328 414
rect 406 397 423 414
rect 447 397 464 414
rect 542 397 559 414
rect 23 151 40 168
rect 195 151 212 168
rect 321 151 338 168
rect 535 149 552 166
rect 10 -40 27 -23
rect 110 -40 127 -23
rect 184 -40 201 -23
rect 281 -40 298 -23
rect 316 -40 333 -23
rect 417 -40 434 -23
rect 452 -40 469 -23
rect 553 -40 570 -23
<< metal1 >>
rect -2 414 577 422
rect -2 397 5 414
rect 22 397 100 414
rect 117 397 175 414
rect 192 397 270 414
rect 287 397 311 414
rect 328 397 406 414
rect 423 397 447 414
rect 464 397 542 414
rect 559 397 577 414
rect -2 389 577 397
rect 17 168 344 174
rect 17 151 23 168
rect 40 151 195 168
rect 212 151 321 168
rect 338 151 344 168
rect 17 145 344 151
rect 529 166 558 172
rect 529 149 535 166
rect 552 149 558 166
rect 529 142 558 149
rect -3 -23 577 -15
rect -3 -40 10 -23
rect 27 -40 110 -23
rect 127 -40 184 -23
rect 201 -40 281 -23
rect 298 -40 316 -23
rect 333 -40 417 -23
rect 434 -40 452 -23
rect 469 -40 553 -23
rect 570 -40 577 -23
rect -3 -48 577 -40
<< comment >>
rect -29 -52 577 452
<< labels >>
flabel metal1 s 139 400 169 415 0 FreeSans 400 0 0 0 vdd
port 0 nsew
flabel metal1 s 273 -44 309 -25 0 FreeSans 400 0 0 0 gnd
port 1 nsew
flabel locali s -19 90 -11 101 0 FreeSans 240 0 0 0 blb
port 2 nsew
flabel locali s 146 90 154 101 0 FreeSans 240 0 0 0 bl
port 3 nsew
flabel locali s 458 84 466 95 0 FreeSans 240 0 0 0 rd_en
port 4 nsew
flabel locali s 108 187 116 198 0 FreeSans 200 0 0 0 net1
flabel locali s 199 155 207 166 0 FreeSans 200 0 0 0 net2
flabel locali s 327 200 335 211 0 FreeSans 200 0 0 0 net3
flabel locali s 538 154 546 160 0 FreeSans 240 0 0 0 dout
port 6 nsew
<< end >>
