6-Transistor SRAM Cell Write Operation

.lib "./libs/models/sky130.lib.spice" tt

*** Inverter 1
XM1 q qbar gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.21
XM2 q qbar vdd vdd sky130_fd_pr__pfet_01v8 w=0.84 l=0.21

*** Inverter 2 
XM3 qbar q gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.21
XM4 qbar q vdd vdd sky130_fd_pr__pfet_01v8 w=0.84 l=0.21

*** Access Transistors
XM5 bl wl q gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.21
XM6 blbar wl qbar gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.21

V1 vdd gnd dc 1.8V

Vwl wl gnd pulse 0 1.8 0 60ps 60ps 20ns 40ns
Vbl bl gnd pulse 0 1.8 0 60ps 60ps 5ns 10ns
Vblbar blbar gnd pulse 1.8 0 0 60ps 60ps 5ns 10ns

.tran 0.1n 100n 
.control
run
plot V(wl)+8 V(bl)+6 V(blbar)+4 V(q)+2 V(qbar)
.endc
.end


