* SKY130 Spice File.
.option scale=1.0u
.include "parameters/lod.spice"
.param
+ lv_dlc_rotweak = .00e-9
+ lvhvt_dlc_rotweak = .00e-9
+ lvt_dlc_rotweak = .00e-9
+ hv_dlc_rotweak = .00e-9
+ sky130_fd_pr__nfet_01v8__dlc_rotweak = lv_dlc_rotweak
+ sky130_fd_pr__esd_nfet_01v8__dlc_rotweak = lv_dlc_rotweak
+ sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak = lvt_dlc_rotweak
+ sky130_fd_pr__pfet_01v8__dlc_rotweak = lv_dlc_rotweak
+ sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak = lvt_dlc_rotweak
+ sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak = lvhvt_dlc_rotweak
+ sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_rotweak = hv_dlc_rotweak
+ sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_rotweak = hv_dlc_rotweak
+ sky130_fd_pr__nfet_03v3_nvt__dlc_rotweak = hv_dlc_rotweak
+ sky130_fd_pr__nfet_05v0_nvt__dlc_rotweak = hv_dlc_rotweak
+ sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak = hv_dlc_rotweak
+ sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak = hv_dlc_rotweak
+ sky130_fd_pr__pfet_g5v0d16v0__dlc_rotweak = hv_dlc_rotweak
+ sky130_fd_pr__special_nfet_pass__dlc_rotweak = lv_dlc_rotweak
+ sky130_fd_pr__special_nfet_pass_lowleakage__dlc_rotweak = lv_dlc_rotweak
+ sky130_fd_pr__special_nfet_pass_flash__dlc_rotweak = hv_dlc_rotweak
+ sky130_fd_pr__special_nfet_latch__dlc_rotweak = lv_dlc_rotweak
+ sky130_fd_pr__special_nfet_latch_lowleakage__dlc_rotweak = lv_dlc_rotweak
+ sky130_fd_pr__special_pfet_pass__dlc_rotweak = lv_dlc_rotweak
+ sky130_fd_pr__special_pfet_pass_lowleakage__dlc_rotweak = lv_dlc_rotweak
+ sky130_fd_bs_flash__special_sonosfet_star__dlc_rotweak = hv_dlc_rotweak
+ sky130_fd_bs_flash__special_sonosfet_original__dlc_rotweak = hv_dlc_rotweak
+ sonos_eeol_dlc_rotweak = hv_dlc_rotweak
+ sonos_peol_dlc_rotweak = hv_dlc_rotweak







