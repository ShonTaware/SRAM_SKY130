magic
tech sky130A
timestamp 1616071127
<< nwell >>
rect 0 382 260 554
<< nmos >>
rect 53 159 68 285
rect 195 159 210 285
rect 76 110 118 125
rect 145 110 187 125
<< pmos >>
rect 53 400 68 455
rect 186 405 201 460
<< ndiff >>
rect 18 277 53 285
rect 18 260 26 277
rect 43 260 53 277
rect 18 184 53 260
rect 18 167 26 184
rect 43 167 53 184
rect 18 159 53 167
rect 68 277 118 285
rect 68 260 93 277
rect 110 260 118 277
rect 68 184 118 260
rect 68 167 93 184
rect 110 167 118 184
rect 68 159 118 167
rect 76 125 118 159
rect 145 277 195 285
rect 145 260 153 277
rect 170 260 195 277
rect 145 184 195 260
rect 145 167 153 184
rect 170 167 195 184
rect 145 159 195 167
rect 210 277 245 285
rect 210 260 220 277
rect 237 260 245 277
rect 210 184 245 260
rect 210 167 220 184
rect 237 167 245 184
rect 210 159 245 167
rect 145 125 187 159
rect 76 100 118 110
rect 76 83 93 100
rect 110 83 118 100
rect 76 76 118 83
rect 145 101 187 110
rect 145 84 153 101
rect 170 84 187 101
rect 145 76 187 84
<< pdiff >>
rect 18 447 53 455
rect 18 430 26 447
rect 43 430 53 447
rect 18 400 53 430
rect 68 425 103 455
rect 68 408 78 425
rect 95 408 103 425
rect 68 400 103 408
rect 151 452 186 460
rect 151 435 159 452
rect 176 435 186 452
rect 151 405 186 435
rect 201 430 236 460
rect 201 413 211 430
rect 228 413 236 430
rect 201 405 236 413
<< ndiffc >>
rect 26 260 43 277
rect 26 167 43 184
rect 93 260 110 277
rect 93 167 110 184
rect 153 260 170 277
rect 153 167 170 184
rect 220 260 237 277
rect 220 167 237 184
rect 93 83 110 100
rect 153 84 170 101
<< pdiffc >>
rect 26 430 43 447
rect 78 408 95 425
rect 159 435 176 452
rect 211 413 228 430
<< psubdiff >>
rect 173 9 214 21
rect 173 -8 185 9
rect 202 -8 214 9
rect 173 -20 214 -8
<< nsubdiff >>
rect 18 517 71 535
rect 18 500 36 517
rect 53 500 71 517
rect 18 482 71 500
<< psubdiffcont >>
rect 185 -8 202 9
<< nsubdiffcont >>
rect 36 500 53 517
<< poly >>
rect 53 455 68 468
rect 186 460 201 473
rect 53 389 68 400
rect 53 381 165 389
rect 53 374 140 381
rect 53 285 68 374
rect 132 364 140 374
rect 157 364 165 381
rect 132 356 165 364
rect 90 327 123 335
rect 90 310 98 327
rect 115 324 123 327
rect 186 324 201 405
rect 115 310 210 324
rect 90 309 210 310
rect 90 302 123 309
rect 195 285 210 309
rect 53 146 68 159
rect 195 146 210 159
rect 0 117 76 125
rect 0 110 26 117
rect 18 100 26 110
rect 43 110 76 117
rect 118 110 145 125
rect 187 110 260 125
rect 43 100 51 110
rect 18 92 51 100
<< polycont >>
rect 140 364 157 381
rect 98 310 115 327
rect 26 100 43 117
<< locali >>
rect 28 521 61 525
rect 0 517 260 521
rect 0 500 36 517
rect 53 500 114 517
rect 131 500 161 517
rect 178 500 211 517
rect 228 500 260 517
rect 0 496 260 500
rect 28 492 61 496
rect 28 455 45 492
rect 18 447 51 455
rect 18 430 26 447
rect 43 430 51 447
rect 151 452 184 460
rect 151 435 159 452
rect 176 435 184 452
rect 211 438 228 496
rect 18 422 51 430
rect 70 425 103 433
rect 70 408 78 425
rect 95 408 103 425
rect 70 400 103 408
rect 151 427 184 435
rect 203 430 236 438
rect 85 335 102 400
rect 151 389 168 427
rect 203 413 211 430
rect 228 413 236 430
rect 203 405 236 413
rect 132 381 168 389
rect 132 364 140 381
rect 157 364 168 381
rect 132 356 168 364
rect 85 327 123 335
rect 85 310 98 327
rect 115 310 123 327
rect 85 302 123 310
rect 85 285 102 302
rect 151 285 168 356
rect 18 277 51 285
rect 18 260 26 277
rect 43 260 51 277
rect 18 231 51 260
rect 85 277 118 285
rect 85 260 93 277
rect 110 260 118 277
rect 85 252 118 260
rect 145 277 178 285
rect 145 260 153 277
rect 170 260 178 277
rect 145 252 178 260
rect 212 277 245 285
rect 212 260 220 277
rect 237 260 245 277
rect 212 231 245 260
rect 18 214 245 231
rect 18 184 51 214
rect 18 167 26 184
rect 43 167 51 184
rect 18 159 51 167
rect 85 184 118 192
rect 85 167 93 184
rect 110 167 118 184
rect 85 159 118 167
rect 145 184 178 192
rect 145 167 153 184
rect 170 167 178 184
rect 145 159 178 167
rect 212 184 245 214
rect 212 167 220 184
rect 237 167 245 184
rect 212 159 245 167
rect 18 117 51 125
rect 18 100 26 117
rect 43 100 51 117
rect 18 92 51 100
rect 85 100 118 108
rect 85 83 93 100
rect 110 83 118 100
rect 85 76 118 83
rect 145 101 178 109
rect 145 84 153 101
rect 170 84 178 101
rect 145 76 178 84
rect 94 69 111 76
rect 145 69 162 76
rect 177 13 210 17
rect 228 13 245 159
rect 0 9 260 13
rect 0 -8 21 9
rect 38 -8 114 9
rect 131 -8 185 9
rect 202 -8 260 9
rect 0 -12 260 -8
rect 177 -16 210 -12
<< viali >>
rect 36 500 53 517
rect 114 500 131 517
rect 161 500 178 517
rect 211 500 228 517
rect 140 364 157 381
rect 98 310 115 327
rect 26 100 43 117
rect 94 52 111 69
rect 145 52 162 69
rect 21 -8 38 9
rect 114 -8 131 9
rect 185 -8 202 9
<< metal1 >>
rect 0 517 260 530
rect 0 500 36 517
rect 53 500 114 517
rect 131 500 161 517
rect 178 500 211 517
rect 228 500 260 517
rect 0 485 260 500
rect 134 381 163 387
rect 134 364 140 381
rect 157 364 163 381
rect 134 358 163 364
rect 92 327 121 333
rect 92 310 98 327
rect 115 310 121 327
rect 92 304 121 310
rect 20 117 49 123
rect 20 107 26 117
rect 18 100 26 107
rect 43 107 49 117
rect 43 100 51 107
rect 18 92 51 100
rect 86 69 118 76
rect 86 52 94 69
rect 111 52 118 69
rect 86 44 118 52
rect 137 69 169 76
rect 137 52 145 69
rect 162 52 169 69
rect 137 44 169 52
rect 0 9 260 21
rect 0 -8 21 9
rect 38 -8 114 9
rect 131 -8 185 9
rect 202 -8 260 9
rect 0 -20 260 -8
<< metal2 >>
rect 53 65 67 554
rect 86 65 118 76
rect 53 51 118 65
rect 53 -20 67 51
rect 86 44 118 51
rect 137 66 169 76
rect 195 66 209 554
rect 137 52 209 66
rect 137 44 169 52
rect 195 -20 209 52
<< labels >>
flabel metal1 s 38 503 49 514 0 FreeSans 200 0 0 0 vdd
port 1 nsew
flabel locali s 143 367 154 378 0 FreeSans 200 0 0 0 qb
port 10 nsew
flabel metal2 s 147 52 158 63 0 FreeSans 200 0 0 0 br
port 16 nsew
flabel metal2 s 89 47 115 73 0 FreeSans 200 0 0 0 bl
port 17 nsew
flabel metal1 s 28 102 39 113 0 FreeSans 200 0 0 0 wl
port 5 nsew
flabel metal1 s 187 -5 198 6 0 FreeSans 200 0 0 0 gnd
port 3 nsew
flabel locali s 102 314 113 325 0 FreeSans 200 0 0 0 q
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 260 509
<< end >>
