VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_2_16_sky130A
   CLASS BLOCK ;
   SIZE 65.08 BY 121.62 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  11.22 -10.1 11.74 -9.58 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  21.88 -10.1 22.4 -9.58 ;
      END
   END din0[1]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -14.2 121.1 -13.68 121.62 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -11.74 121.1 -11.22 121.62 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -13.38 121.1 -12.86 121.62 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -12.56 121.1 -12.04 121.62 ;
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  -56.84 -7.64 -56.32 -7.12 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  -56.84 -4.36 -56.32 -3.84 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -25.68 -10.1 -25.16 -9.58 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m3 ;
         RECT  64.52 9.58 65.04 10.1 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m3 ;
         RECT  64.52 11.22 65.04 11.74 ;
      END
   END dout0[1]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  -56.84 -6.0 -55.5 -4.66 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  -56.84 -10.1 -55.5 -8.76 ;
      END
   END gnd
   OBS
   LAYER  m1 ;
      RECT  49.57 37.39 49.86 37.68 ;
      RECT  50.02 34.79 50.34 35.11 ;
      RECT  48.83 35.27 49.16 35.42 ;
      RECT  48.65 34.15 51.25 34.56 ;
      RECT  48.65 39.2 51.25 39.65 ;
      RECT  49.51 34.79 49.83 35.11 ;
      RECT  49.99 37.93 50.28 38.22 ;
      RECT  48.85 35.42 49.14 35.58 ;
      RECT  49.57 41.49 49.86 41.2 ;
      RECT  50.02 44.09 50.34 43.77 ;
      RECT  48.83 43.61 49.16 43.46 ;
      RECT  48.65 44.73 51.25 44.32 ;
      RECT  48.65 39.68 51.25 39.23 ;
      RECT  49.51 44.09 49.83 43.77 ;
      RECT  49.99 40.95 50.28 40.66 ;
      RECT  48.85 43.46 49.14 43.3 ;
      RECT  49.57 47.57 49.86 47.86 ;
      RECT  50.02 44.97 50.34 45.29 ;
      RECT  48.83 45.45 49.16 45.6 ;
      RECT  48.65 44.33 51.25 44.74 ;
      RECT  48.65 49.38 51.25 49.83 ;
      RECT  49.51 44.97 49.83 45.29 ;
      RECT  49.99 48.11 50.28 48.4 ;
      RECT  48.85 45.6 49.14 45.76 ;
      RECT  49.57 51.67 49.86 51.38 ;
      RECT  50.02 54.27 50.34 53.95 ;
      RECT  48.83 53.79 49.16 53.64 ;
      RECT  48.65 54.91 51.25 54.5 ;
      RECT  48.65 49.86 51.25 49.41 ;
      RECT  49.51 54.27 49.83 53.95 ;
      RECT  49.99 51.13 50.28 50.84 ;
      RECT  48.85 53.64 49.14 53.48 ;
      RECT  49.57 57.75 49.86 58.04 ;
      RECT  50.02 55.15 50.34 55.47 ;
      RECT  48.83 55.63 49.16 55.78 ;
      RECT  48.65 54.51 51.25 54.92 ;
      RECT  48.65 59.56 51.25 60.01 ;
      RECT  49.51 55.15 49.83 55.47 ;
      RECT  49.99 58.29 50.28 58.58 ;
      RECT  48.85 55.78 49.14 55.94 ;
      RECT  49.57 61.85 49.86 61.56 ;
      RECT  50.02 64.45 50.34 64.13 ;
      RECT  48.83 63.97 49.16 63.82 ;
      RECT  48.65 65.09 51.25 64.68 ;
      RECT  48.65 60.04 51.25 59.59 ;
      RECT  49.51 64.45 49.83 64.13 ;
      RECT  49.99 61.31 50.28 61.02 ;
      RECT  48.85 63.82 49.14 63.66 ;
      RECT  49.57 67.93 49.86 68.22 ;
      RECT  50.02 65.33 50.34 65.65 ;
      RECT  48.83 65.81 49.16 65.96 ;
      RECT  48.65 64.69 51.25 65.1 ;
      RECT  48.65 69.74 51.25 70.19 ;
      RECT  49.51 65.33 49.83 65.65 ;
      RECT  49.99 68.47 50.28 68.76 ;
      RECT  48.85 65.96 49.14 66.12 ;
      RECT  49.57 72.03 49.86 71.74 ;
      RECT  50.02 74.63 50.34 74.31 ;
      RECT  48.83 74.15 49.16 74.0 ;
      RECT  48.65 75.27 51.25 74.86 ;
      RECT  48.65 70.22 51.25 69.77 ;
      RECT  49.51 74.63 49.83 74.31 ;
      RECT  49.99 71.49 50.28 71.2 ;
      RECT  48.85 74.0 49.14 73.84 ;
      RECT  49.57 78.11 49.86 78.4 ;
      RECT  50.02 75.51 50.34 75.83 ;
      RECT  48.83 75.99 49.16 76.14 ;
      RECT  48.65 74.87 51.25 75.28 ;
      RECT  48.65 79.92 51.25 80.37 ;
      RECT  49.51 75.51 49.83 75.83 ;
      RECT  49.99 78.65 50.28 78.94 ;
      RECT  48.85 76.14 49.14 76.3 ;
      RECT  49.57 82.21 49.86 81.92 ;
      RECT  50.02 84.81 50.34 84.49 ;
      RECT  48.83 84.33 49.16 84.18 ;
      RECT  48.65 85.45 51.25 85.04 ;
      RECT  48.65 80.4 51.25 79.95 ;
      RECT  49.51 84.81 49.83 84.49 ;
      RECT  49.99 81.67 50.28 81.38 ;
      RECT  48.85 84.18 49.14 84.02 ;
      RECT  49.57 88.29 49.86 88.58 ;
      RECT  50.02 85.69 50.34 86.01 ;
      RECT  48.83 86.17 49.16 86.32 ;
      RECT  48.65 85.05 51.25 85.46 ;
      RECT  48.65 90.1 51.25 90.55 ;
      RECT  49.51 85.69 49.83 86.01 ;
      RECT  49.99 88.83 50.28 89.12 ;
      RECT  48.85 86.32 49.14 86.48 ;
      RECT  49.57 92.39 49.86 92.1 ;
      RECT  50.02 94.99 50.34 94.67 ;
      RECT  48.83 94.51 49.16 94.36 ;
      RECT  48.65 95.63 51.25 95.22 ;
      RECT  48.65 90.58 51.25 90.13 ;
      RECT  49.51 94.99 49.83 94.67 ;
      RECT  49.99 91.85 50.28 91.56 ;
      RECT  48.85 94.36 49.14 94.2 ;
      RECT  49.57 98.47 49.86 98.76 ;
      RECT  50.02 95.87 50.34 96.19 ;
      RECT  48.83 96.35 49.16 96.5 ;
      RECT  48.65 95.23 51.25 95.64 ;
      RECT  48.65 100.28 51.25 100.73 ;
      RECT  49.51 95.87 49.83 96.19 ;
      RECT  49.99 99.01 50.28 99.3 ;
      RECT  48.85 96.5 49.14 96.66 ;
      RECT  49.57 102.57 49.86 102.28 ;
      RECT  50.02 105.17 50.34 104.85 ;
      RECT  48.83 104.69 49.16 104.54 ;
      RECT  48.65 105.81 51.25 105.4 ;
      RECT  48.65 100.76 51.25 100.31 ;
      RECT  49.51 105.17 49.83 104.85 ;
      RECT  49.99 102.03 50.28 101.74 ;
      RECT  48.85 104.54 49.14 104.38 ;
      RECT  49.57 108.65 49.86 108.94 ;
      RECT  50.02 106.05 50.34 106.37 ;
      RECT  48.83 106.53 49.16 106.68 ;
      RECT  48.65 105.41 51.25 105.82 ;
      RECT  48.65 110.46 51.25 110.91 ;
      RECT  49.51 106.05 49.83 106.37 ;
      RECT  49.99 109.19 50.28 109.48 ;
      RECT  48.85 106.68 49.14 106.84 ;
      RECT  49.57 112.75 49.86 112.46 ;
      RECT  50.02 115.35 50.34 115.03 ;
      RECT  48.83 114.87 49.16 114.72 ;
      RECT  48.65 115.99 51.25 115.58 ;
      RECT  48.65 110.94 51.25 110.49 ;
      RECT  49.51 115.35 49.83 115.03 ;
      RECT  49.99 112.21 50.28 111.92 ;
      RECT  48.85 114.72 49.14 114.56 ;
      RECT  52.17 37.39 52.46 37.68 ;
      RECT  52.62 34.79 52.94 35.11 ;
      RECT  51.43 35.27 51.76 35.42 ;
      RECT  51.25 34.15 53.85 34.56 ;
      RECT  51.25 39.2 53.85 39.65 ;
      RECT  52.11 34.79 52.43 35.11 ;
      RECT  52.59 37.93 52.88 38.22 ;
      RECT  51.45 35.42 51.74 35.58 ;
      RECT  52.17 41.49 52.46 41.2 ;
      RECT  52.62 44.09 52.94 43.77 ;
      RECT  51.43 43.61 51.76 43.46 ;
      RECT  51.25 44.73 53.85 44.32 ;
      RECT  51.25 39.68 53.85 39.23 ;
      RECT  52.11 44.09 52.43 43.77 ;
      RECT  52.59 40.95 52.88 40.66 ;
      RECT  51.45 43.46 51.74 43.3 ;
      RECT  52.17 47.57 52.46 47.86 ;
      RECT  52.62 44.97 52.94 45.29 ;
      RECT  51.43 45.45 51.76 45.6 ;
      RECT  51.25 44.33 53.85 44.74 ;
      RECT  51.25 49.38 53.85 49.83 ;
      RECT  52.11 44.97 52.43 45.29 ;
      RECT  52.59 48.11 52.88 48.4 ;
      RECT  51.45 45.6 51.74 45.76 ;
      RECT  52.17 51.67 52.46 51.38 ;
      RECT  52.62 54.27 52.94 53.95 ;
      RECT  51.43 53.79 51.76 53.64 ;
      RECT  51.25 54.91 53.85 54.5 ;
      RECT  51.25 49.86 53.85 49.41 ;
      RECT  52.11 54.27 52.43 53.95 ;
      RECT  52.59 51.13 52.88 50.84 ;
      RECT  51.45 53.64 51.74 53.48 ;
      RECT  52.17 57.75 52.46 58.04 ;
      RECT  52.62 55.15 52.94 55.47 ;
      RECT  51.43 55.63 51.76 55.78 ;
      RECT  51.25 54.51 53.85 54.92 ;
      RECT  51.25 59.56 53.85 60.01 ;
      RECT  52.11 55.15 52.43 55.47 ;
      RECT  52.59 58.29 52.88 58.58 ;
      RECT  51.45 55.78 51.74 55.94 ;
      RECT  52.17 61.85 52.46 61.56 ;
      RECT  52.62 64.45 52.94 64.13 ;
      RECT  51.43 63.97 51.76 63.82 ;
      RECT  51.25 65.09 53.85 64.68 ;
      RECT  51.25 60.04 53.85 59.59 ;
      RECT  52.11 64.45 52.43 64.13 ;
      RECT  52.59 61.31 52.88 61.02 ;
      RECT  51.45 63.82 51.74 63.66 ;
      RECT  52.17 67.93 52.46 68.22 ;
      RECT  52.62 65.33 52.94 65.65 ;
      RECT  51.43 65.81 51.76 65.96 ;
      RECT  51.25 64.69 53.85 65.1 ;
      RECT  51.25 69.74 53.85 70.19 ;
      RECT  52.11 65.33 52.43 65.65 ;
      RECT  52.59 68.47 52.88 68.76 ;
      RECT  51.45 65.96 51.74 66.12 ;
      RECT  52.17 72.03 52.46 71.74 ;
      RECT  52.62 74.63 52.94 74.31 ;
      RECT  51.43 74.15 51.76 74.0 ;
      RECT  51.25 75.27 53.85 74.86 ;
      RECT  51.25 70.22 53.85 69.77 ;
      RECT  52.11 74.63 52.43 74.31 ;
      RECT  52.59 71.49 52.88 71.2 ;
      RECT  51.45 74.0 51.74 73.84 ;
      RECT  52.17 78.11 52.46 78.4 ;
      RECT  52.62 75.51 52.94 75.83 ;
      RECT  51.43 75.99 51.76 76.14 ;
      RECT  51.25 74.87 53.85 75.28 ;
      RECT  51.25 79.92 53.85 80.37 ;
      RECT  52.11 75.51 52.43 75.83 ;
      RECT  52.59 78.65 52.88 78.94 ;
      RECT  51.45 76.14 51.74 76.3 ;
      RECT  52.17 82.21 52.46 81.92 ;
      RECT  52.62 84.81 52.94 84.49 ;
      RECT  51.43 84.33 51.76 84.18 ;
      RECT  51.25 85.45 53.85 85.04 ;
      RECT  51.25 80.4 53.85 79.95 ;
      RECT  52.11 84.81 52.43 84.49 ;
      RECT  52.59 81.67 52.88 81.38 ;
      RECT  51.45 84.18 51.74 84.02 ;
      RECT  52.17 88.29 52.46 88.58 ;
      RECT  52.62 85.69 52.94 86.01 ;
      RECT  51.43 86.17 51.76 86.32 ;
      RECT  51.25 85.05 53.85 85.46 ;
      RECT  51.25 90.1 53.85 90.55 ;
      RECT  52.11 85.69 52.43 86.01 ;
      RECT  52.59 88.83 52.88 89.12 ;
      RECT  51.45 86.32 51.74 86.48 ;
      RECT  52.17 92.39 52.46 92.1 ;
      RECT  52.62 94.99 52.94 94.67 ;
      RECT  51.43 94.51 51.76 94.36 ;
      RECT  51.25 95.63 53.85 95.22 ;
      RECT  51.25 90.58 53.85 90.13 ;
      RECT  52.11 94.99 52.43 94.67 ;
      RECT  52.59 91.85 52.88 91.56 ;
      RECT  51.45 94.36 51.74 94.2 ;
      RECT  52.17 98.47 52.46 98.76 ;
      RECT  52.62 95.87 52.94 96.19 ;
      RECT  51.43 96.35 51.76 96.5 ;
      RECT  51.25 95.23 53.85 95.64 ;
      RECT  51.25 100.28 53.85 100.73 ;
      RECT  52.11 95.87 52.43 96.19 ;
      RECT  52.59 99.01 52.88 99.3 ;
      RECT  51.45 96.5 51.74 96.66 ;
      RECT  52.17 102.57 52.46 102.28 ;
      RECT  52.62 105.17 52.94 104.85 ;
      RECT  51.43 104.69 51.76 104.54 ;
      RECT  51.25 105.81 53.85 105.4 ;
      RECT  51.25 100.76 53.85 100.31 ;
      RECT  52.11 105.17 52.43 104.85 ;
      RECT  52.59 102.03 52.88 101.74 ;
      RECT  51.45 104.54 51.74 104.38 ;
      RECT  52.17 108.65 52.46 108.94 ;
      RECT  52.62 106.05 52.94 106.37 ;
      RECT  51.43 106.53 51.76 106.68 ;
      RECT  51.25 105.41 53.85 105.82 ;
      RECT  51.25 110.46 53.85 110.91 ;
      RECT  52.11 106.05 52.43 106.37 ;
      RECT  52.59 109.19 52.88 109.48 ;
      RECT  51.45 106.68 51.74 106.84 ;
      RECT  52.17 112.75 52.46 112.46 ;
      RECT  52.62 115.35 52.94 115.03 ;
      RECT  51.43 114.87 51.76 114.72 ;
      RECT  51.25 115.99 53.85 115.58 ;
      RECT  51.25 110.94 53.85 110.49 ;
      RECT  52.11 115.35 52.43 115.03 ;
      RECT  52.59 112.21 52.88 111.92 ;
      RECT  51.45 114.72 51.74 114.56 ;
      RECT  48.65 35.42 53.85 35.58 ;
      RECT  48.65 43.3 53.85 43.46 ;
      RECT  48.65 45.6 53.85 45.76 ;
      RECT  48.65 53.48 53.85 53.64 ;
      RECT  48.65 55.78 53.85 55.94 ;
      RECT  48.65 63.66 53.85 63.82 ;
      RECT  48.65 65.96 53.85 66.12 ;
      RECT  48.65 73.84 53.85 74.0 ;
      RECT  48.65 76.14 53.85 76.3 ;
      RECT  48.65 84.02 53.85 84.18 ;
      RECT  48.65 86.32 53.85 86.48 ;
      RECT  48.65 94.2 53.85 94.36 ;
      RECT  48.65 96.5 53.85 96.66 ;
      RECT  48.65 104.38 53.85 104.54 ;
      RECT  48.65 106.68 53.85 106.84 ;
      RECT  48.65 114.56 53.85 114.72 ;
      RECT  51.25 79.92 53.85 80.37 ;
      RECT  48.65 100.31 51.25 100.76 ;
      RECT  48.65 79.95 51.25 80.4 ;
      RECT  51.25 39.2 53.85 39.65 ;
      RECT  48.65 49.38 51.25 49.83 ;
      RECT  48.65 69.74 51.25 70.19 ;
      RECT  51.25 69.77 53.85 70.22 ;
      RECT  48.65 110.46 51.25 110.91 ;
      RECT  51.25 69.74 53.85 70.19 ;
      RECT  48.65 79.92 51.25 80.37 ;
      RECT  51.25 49.41 53.85 49.86 ;
      RECT  51.25 79.95 53.85 80.4 ;
      RECT  48.65 69.77 51.25 70.22 ;
      RECT  51.25 90.1 53.85 90.55 ;
      RECT  51.25 110.49 53.85 110.94 ;
      RECT  51.25 110.46 53.85 110.91 ;
      RECT  48.65 39.2 51.25 39.65 ;
      RECT  51.25 90.13 53.85 90.58 ;
      RECT  48.65 110.49 51.25 110.94 ;
      RECT  51.25 100.31 53.85 100.76 ;
      RECT  48.65 90.13 51.25 90.58 ;
      RECT  51.25 49.38 53.85 49.83 ;
      RECT  48.65 49.41 51.25 49.86 ;
      RECT  48.65 39.23 51.25 39.68 ;
      RECT  51.25 39.23 53.85 39.68 ;
      RECT  48.65 90.1 51.25 90.55 ;
      RECT  48.65 59.56 51.25 60.01 ;
      RECT  48.65 59.59 51.25 60.04 ;
      RECT  51.25 59.59 53.85 60.04 ;
      RECT  51.25 59.56 53.85 60.01 ;
      RECT  51.25 100.28 53.85 100.73 ;
      RECT  48.65 100.28 51.25 100.73 ;
      RECT  51.25 44.33 53.85 44.74 ;
      RECT  51.25 85.04 53.85 85.45 ;
      RECT  48.65 105.4 51.25 105.81 ;
      RECT  48.65 44.32 51.25 44.73 ;
      RECT  51.25 74.87 53.85 75.28 ;
      RECT  48.65 54.5 51.25 54.91 ;
      RECT  51.25 105.4 53.85 105.81 ;
      RECT  51.25 115.58 53.85 115.99 ;
      RECT  48.65 74.87 51.25 75.28 ;
      RECT  51.25 95.23 53.85 95.64 ;
      RECT  48.65 74.86 51.25 75.27 ;
      RECT  48.65 105.41 51.25 105.82 ;
      RECT  48.65 85.05 51.25 85.46 ;
      RECT  51.25 105.41 53.85 105.82 ;
      RECT  48.65 95.23 51.25 95.64 ;
      RECT  51.25 95.22 53.85 95.63 ;
      RECT  51.25 64.68 53.85 65.09 ;
      RECT  48.65 115.58 51.25 115.99 ;
      RECT  48.65 44.33 51.25 44.74 ;
      RECT  51.25 74.86 53.85 75.27 ;
      RECT  48.65 64.68 51.25 65.09 ;
      RECT  48.65 64.69 51.25 65.1 ;
      RECT  48.65 34.15 51.25 34.56 ;
      RECT  51.25 34.15 53.85 34.56 ;
      RECT  51.25 44.32 53.85 44.73 ;
      RECT  48.65 85.04 51.25 85.45 ;
      RECT  51.25 85.05 53.85 85.46 ;
      RECT  48.65 95.22 51.25 95.63 ;
      RECT  51.25 64.69 53.85 65.1 ;
      RECT  48.65 54.51 51.25 54.92 ;
      RECT  51.25 54.51 53.85 54.92 ;
      RECT  51.25 54.5 53.85 54.91 ;
      RECT  46.97 27.21 47.26 27.5 ;
      RECT  47.42 24.61 47.74 24.93 ;
      RECT  46.23 25.09 46.56 25.24 ;
      RECT  46.05 23.97 48.65 24.38 ;
      RECT  46.05 29.02 48.65 29.47 ;
      RECT  46.91 24.61 47.23 24.93 ;
      RECT  47.39 27.75 47.68 28.04 ;
      RECT  46.25 25.24 46.54 25.4 ;
      RECT  46.97 31.31 47.26 31.02 ;
      RECT  47.42 33.91 47.74 33.59 ;
      RECT  46.23 33.43 46.56 33.28 ;
      RECT  46.05 34.55 48.65 34.14 ;
      RECT  46.05 29.5 48.65 29.05 ;
      RECT  46.91 33.91 47.23 33.59 ;
      RECT  47.39 30.77 47.68 30.48 ;
      RECT  46.25 33.28 46.54 33.12 ;
      RECT  46.97 37.39 47.26 37.68 ;
      RECT  47.42 34.79 47.74 35.11 ;
      RECT  46.23 35.27 46.56 35.42 ;
      RECT  46.05 34.15 48.65 34.56 ;
      RECT  46.05 39.2 48.65 39.65 ;
      RECT  46.91 34.79 47.23 35.11 ;
      RECT  47.39 37.93 47.68 38.22 ;
      RECT  46.25 35.42 46.54 35.58 ;
      RECT  46.97 41.49 47.26 41.2 ;
      RECT  47.42 44.09 47.74 43.77 ;
      RECT  46.23 43.61 46.56 43.46 ;
      RECT  46.05 44.73 48.65 44.32 ;
      RECT  46.05 39.68 48.65 39.23 ;
      RECT  46.91 44.09 47.23 43.77 ;
      RECT  47.39 40.95 47.68 40.66 ;
      RECT  46.25 43.46 46.54 43.3 ;
      RECT  46.97 47.57 47.26 47.86 ;
      RECT  47.42 44.97 47.74 45.29 ;
      RECT  46.23 45.45 46.56 45.6 ;
      RECT  46.05 44.33 48.65 44.74 ;
      RECT  46.05 49.38 48.65 49.83 ;
      RECT  46.91 44.97 47.23 45.29 ;
      RECT  47.39 48.11 47.68 48.4 ;
      RECT  46.25 45.6 46.54 45.76 ;
      RECT  46.97 51.67 47.26 51.38 ;
      RECT  47.42 54.27 47.74 53.95 ;
      RECT  46.23 53.79 46.56 53.64 ;
      RECT  46.05 54.91 48.65 54.5 ;
      RECT  46.05 49.86 48.65 49.41 ;
      RECT  46.91 54.27 47.23 53.95 ;
      RECT  47.39 51.13 47.68 50.84 ;
      RECT  46.25 53.64 46.54 53.48 ;
      RECT  46.97 57.75 47.26 58.04 ;
      RECT  47.42 55.15 47.74 55.47 ;
      RECT  46.23 55.63 46.56 55.78 ;
      RECT  46.05 54.51 48.65 54.92 ;
      RECT  46.05 59.56 48.65 60.01 ;
      RECT  46.91 55.15 47.23 55.47 ;
      RECT  47.39 58.29 47.68 58.58 ;
      RECT  46.25 55.78 46.54 55.94 ;
      RECT  46.97 61.85 47.26 61.56 ;
      RECT  47.42 64.45 47.74 64.13 ;
      RECT  46.23 63.97 46.56 63.82 ;
      RECT  46.05 65.09 48.65 64.68 ;
      RECT  46.05 60.04 48.65 59.59 ;
      RECT  46.91 64.45 47.23 64.13 ;
      RECT  47.39 61.31 47.68 61.02 ;
      RECT  46.25 63.82 46.54 63.66 ;
      RECT  46.97 67.93 47.26 68.22 ;
      RECT  47.42 65.33 47.74 65.65 ;
      RECT  46.23 65.81 46.56 65.96 ;
      RECT  46.05 64.69 48.65 65.1 ;
      RECT  46.05 69.74 48.65 70.19 ;
      RECT  46.91 65.33 47.23 65.65 ;
      RECT  47.39 68.47 47.68 68.76 ;
      RECT  46.25 65.96 46.54 66.12 ;
      RECT  46.97 72.03 47.26 71.74 ;
      RECT  47.42 74.63 47.74 74.31 ;
      RECT  46.23 74.15 46.56 74.0 ;
      RECT  46.05 75.27 48.65 74.86 ;
      RECT  46.05 70.22 48.65 69.77 ;
      RECT  46.91 74.63 47.23 74.31 ;
      RECT  47.39 71.49 47.68 71.2 ;
      RECT  46.25 74.0 46.54 73.84 ;
      RECT  46.97 78.11 47.26 78.4 ;
      RECT  47.42 75.51 47.74 75.83 ;
      RECT  46.23 75.99 46.56 76.14 ;
      RECT  46.05 74.87 48.65 75.28 ;
      RECT  46.05 79.92 48.65 80.37 ;
      RECT  46.91 75.51 47.23 75.83 ;
      RECT  47.39 78.65 47.68 78.94 ;
      RECT  46.25 76.14 46.54 76.3 ;
      RECT  46.97 82.21 47.26 81.92 ;
      RECT  47.42 84.81 47.74 84.49 ;
      RECT  46.23 84.33 46.56 84.18 ;
      RECT  46.05 85.45 48.65 85.04 ;
      RECT  46.05 80.4 48.65 79.95 ;
      RECT  46.91 84.81 47.23 84.49 ;
      RECT  47.39 81.67 47.68 81.38 ;
      RECT  46.25 84.18 46.54 84.02 ;
      RECT  46.97 88.29 47.26 88.58 ;
      RECT  47.42 85.69 47.74 86.01 ;
      RECT  46.23 86.17 46.56 86.32 ;
      RECT  46.05 85.05 48.65 85.46 ;
      RECT  46.05 90.1 48.65 90.55 ;
      RECT  46.91 85.69 47.23 86.01 ;
      RECT  47.39 88.83 47.68 89.12 ;
      RECT  46.25 86.32 46.54 86.48 ;
      RECT  46.97 92.39 47.26 92.1 ;
      RECT  47.42 94.99 47.74 94.67 ;
      RECT  46.23 94.51 46.56 94.36 ;
      RECT  46.05 95.63 48.65 95.22 ;
      RECT  46.05 90.58 48.65 90.13 ;
      RECT  46.91 94.99 47.23 94.67 ;
      RECT  47.39 91.85 47.68 91.56 ;
      RECT  46.25 94.36 46.54 94.2 ;
      RECT  46.97 98.47 47.26 98.76 ;
      RECT  47.42 95.87 47.74 96.19 ;
      RECT  46.23 96.35 46.56 96.5 ;
      RECT  46.05 95.23 48.65 95.64 ;
      RECT  46.05 100.28 48.65 100.73 ;
      RECT  46.91 95.87 47.23 96.19 ;
      RECT  47.39 99.01 47.68 99.3 ;
      RECT  46.25 96.5 46.54 96.66 ;
      RECT  46.97 102.57 47.26 102.28 ;
      RECT  47.42 105.17 47.74 104.85 ;
      RECT  46.23 104.69 46.56 104.54 ;
      RECT  46.05 105.81 48.65 105.4 ;
      RECT  46.05 100.76 48.65 100.31 ;
      RECT  46.91 105.17 47.23 104.85 ;
      RECT  47.39 102.03 47.68 101.74 ;
      RECT  46.25 104.54 46.54 104.38 ;
      RECT  46.97 108.65 47.26 108.94 ;
      RECT  47.42 106.05 47.74 106.37 ;
      RECT  46.23 106.53 46.56 106.68 ;
      RECT  46.05 105.41 48.65 105.82 ;
      RECT  46.05 110.46 48.65 110.91 ;
      RECT  46.91 106.05 47.23 106.37 ;
      RECT  47.39 109.19 47.68 109.48 ;
      RECT  46.25 106.68 46.54 106.84 ;
      RECT  46.97 112.75 47.26 112.46 ;
      RECT  47.42 115.35 47.74 115.03 ;
      RECT  46.23 114.87 46.56 114.72 ;
      RECT  46.05 115.99 48.65 115.58 ;
      RECT  46.05 110.94 48.65 110.49 ;
      RECT  46.91 115.35 47.23 115.03 ;
      RECT  47.39 112.21 47.68 111.92 ;
      RECT  46.25 114.72 46.54 114.56 ;
      RECT  46.97 118.83 47.26 119.12 ;
      RECT  47.42 116.23 47.74 116.55 ;
      RECT  46.23 116.71 46.56 116.86 ;
      RECT  46.05 115.59 48.65 116.0 ;
      RECT  46.05 120.64 48.65 121.09 ;
      RECT  46.91 116.23 47.23 116.55 ;
      RECT  47.39 119.37 47.68 119.66 ;
      RECT  46.25 116.86 46.54 117.02 ;
      RECT  46.05 25.24 48.65 25.4 ;
      RECT  46.05 33.12 48.65 33.28 ;
      RECT  46.05 35.42 48.65 35.58 ;
      RECT  46.05 43.3 48.65 43.46 ;
      RECT  46.05 45.6 48.65 45.76 ;
      RECT  46.05 53.48 48.65 53.64 ;
      RECT  46.05 55.78 48.65 55.94 ;
      RECT  46.05 63.66 48.65 63.82 ;
      RECT  46.05 65.96 48.65 66.12 ;
      RECT  46.05 73.84 48.65 74.0 ;
      RECT  46.05 76.14 48.65 76.3 ;
      RECT  46.05 84.02 48.65 84.18 ;
      RECT  46.05 86.32 48.65 86.48 ;
      RECT  46.05 94.2 48.65 94.36 ;
      RECT  46.05 96.5 48.65 96.66 ;
      RECT  46.05 104.38 48.65 104.54 ;
      RECT  46.05 106.68 48.65 106.84 ;
      RECT  46.05 114.56 48.65 114.72 ;
      RECT  46.05 116.86 48.65 117.02 ;
      RECT  46.05 90.13 48.65 90.58 ;
      RECT  46.05 69.77 48.65 70.22 ;
      RECT  46.05 39.2 48.65 39.65 ;
      RECT  46.05 59.56 48.65 60.01 ;
      RECT  46.05 100.28 48.65 100.73 ;
      RECT  46.05 110.49 48.65 110.94 ;
      RECT  46.05 69.74 48.65 70.19 ;
      RECT  46.05 59.59 48.65 60.04 ;
      RECT  46.05 100.31 48.65 100.76 ;
      RECT  46.05 79.95 48.65 80.4 ;
      RECT  46.05 110.46 48.65 110.91 ;
      RECT  46.05 39.23 48.65 39.68 ;
      RECT  46.05 29.05 48.65 29.5 ;
      RECT  46.05 79.92 48.65 80.37 ;
      RECT  46.05 49.38 48.65 49.83 ;
      RECT  46.05 49.41 48.65 49.86 ;
      RECT  46.05 90.1 48.65 90.55 ;
      RECT  46.05 105.41 48.65 105.82 ;
      RECT  46.05 95.22 48.65 95.63 ;
      RECT  46.05 34.14 48.65 34.55 ;
      RECT  46.05 44.32 48.65 44.73 ;
      RECT  46.05 64.69 48.65 65.1 ;
      RECT  46.05 64.68 48.65 65.09 ;
      RECT  46.05 95.23 48.65 95.64 ;
      RECT  46.05 74.87 48.65 75.28 ;
      RECT  46.05 85.05 48.65 85.46 ;
      RECT  46.05 105.4 48.65 105.81 ;
      RECT  46.05 34.15 48.65 34.56 ;
      RECT  46.05 54.5 48.65 54.91 ;
      RECT  46.05 54.51 48.65 54.92 ;
      RECT  46.05 115.58 48.65 115.99 ;
      RECT  46.05 74.86 48.65 75.27 ;
      RECT  46.05 85.04 48.65 85.45 ;
      RECT  46.05 44.33 48.65 44.74 ;
      RECT  49.57 31.31 49.86 31.02 ;
      RECT  50.02 33.91 50.34 33.59 ;
      RECT  48.83 33.43 49.16 33.28 ;
      RECT  48.65 34.55 51.25 34.14 ;
      RECT  48.65 29.5 51.25 29.05 ;
      RECT  49.51 33.91 49.83 33.59 ;
      RECT  49.99 30.77 50.28 30.48 ;
      RECT  48.85 33.28 49.14 33.12 ;
      RECT  52.17 31.31 52.46 31.02 ;
      RECT  52.62 33.91 52.94 33.59 ;
      RECT  51.43 33.43 51.76 33.28 ;
      RECT  51.25 34.55 53.85 34.14 ;
      RECT  51.25 29.5 53.85 29.05 ;
      RECT  52.11 33.91 52.43 33.59 ;
      RECT  52.59 30.77 52.88 30.48 ;
      RECT  51.45 33.28 51.74 33.12 ;
      RECT  48.65 33.28 53.85 33.12 ;
      RECT  51.25 29.5 53.85 29.05 ;
      RECT  48.65 29.5 51.25 29.05 ;
      RECT  48.65 34.55 51.25 34.14 ;
      RECT  51.25 34.55 53.85 34.14 ;
      RECT  49.57 27.21 49.86 27.5 ;
      RECT  50.02 24.61 50.34 24.93 ;
      RECT  48.83 25.09 49.16 25.24 ;
      RECT  48.65 23.97 51.25 24.38 ;
      RECT  48.65 29.02 51.25 29.47 ;
      RECT  49.51 24.61 49.83 24.93 ;
      RECT  49.99 27.75 50.28 28.04 ;
      RECT  48.85 25.24 49.14 25.4 ;
      RECT  52.17 27.21 52.46 27.5 ;
      RECT  52.62 24.61 52.94 24.93 ;
      RECT  51.43 25.09 51.76 25.24 ;
      RECT  51.25 23.97 53.85 24.38 ;
      RECT  51.25 29.02 53.85 29.47 ;
      RECT  52.11 24.61 52.43 24.93 ;
      RECT  52.59 27.75 52.88 28.04 ;
      RECT  51.45 25.24 51.74 25.4 ;
      RECT  48.65 25.24 53.85 25.4 ;
      RECT  51.25 29.02 53.85 29.47 ;
      RECT  48.65 29.02 51.25 29.47 ;
      RECT  48.65 23.97 51.25 24.38 ;
      RECT  51.25 23.97 53.85 24.38 ;
      RECT  49.57 118.83 49.86 119.12 ;
      RECT  50.02 116.23 50.34 116.55 ;
      RECT  48.83 116.71 49.16 116.86 ;
      RECT  48.65 115.59 51.25 116.0 ;
      RECT  48.65 120.64 51.25 121.09 ;
      RECT  49.51 116.23 49.83 116.55 ;
      RECT  49.99 119.37 50.28 119.66 ;
      RECT  48.85 116.86 49.14 117.02 ;
      RECT  52.17 118.83 52.46 119.12 ;
      RECT  52.62 116.23 52.94 116.55 ;
      RECT  51.43 116.71 51.76 116.86 ;
      RECT  51.25 115.59 53.85 116.0 ;
      RECT  51.25 120.64 53.85 121.09 ;
      RECT  52.11 116.23 52.43 116.55 ;
      RECT  52.59 119.37 52.88 119.66 ;
      RECT  51.45 116.86 51.74 117.02 ;
      RECT  48.65 116.86 53.85 117.02 ;
      RECT  51.25 120.64 53.85 121.09 ;
      RECT  48.65 120.64 51.25 121.09 ;
      RECT  48.65 115.59 51.25 116.0 ;
      RECT  51.25 115.59 53.85 116.0 ;
      RECT  44.37 27.21 44.66 27.5 ;
      RECT  44.82 24.61 45.14 24.93 ;
      RECT  43.63 25.09 43.96 25.24 ;
      RECT  43.45 23.97 46.05 24.38 ;
      RECT  43.45 29.02 46.05 29.47 ;
      RECT  44.31 24.61 44.63 24.93 ;
      RECT  44.79 27.75 45.08 28.04 ;
      RECT  43.65 25.24 43.94 25.4 ;
      RECT  44.37 31.31 44.66 31.02 ;
      RECT  44.82 33.91 45.14 33.59 ;
      RECT  43.63 33.43 43.96 33.28 ;
      RECT  43.45 34.55 46.05 34.14 ;
      RECT  43.45 29.5 46.05 29.05 ;
      RECT  44.31 33.91 44.63 33.59 ;
      RECT  44.79 30.77 45.08 30.48 ;
      RECT  43.65 33.28 43.94 33.12 ;
      RECT  44.37 37.39 44.66 37.68 ;
      RECT  44.82 34.79 45.14 35.11 ;
      RECT  43.63 35.27 43.96 35.42 ;
      RECT  43.45 34.15 46.05 34.56 ;
      RECT  43.45 39.2 46.05 39.65 ;
      RECT  44.31 34.79 44.63 35.11 ;
      RECT  44.79 37.93 45.08 38.22 ;
      RECT  43.65 35.42 43.94 35.58 ;
      RECT  44.37 41.49 44.66 41.2 ;
      RECT  44.82 44.09 45.14 43.77 ;
      RECT  43.63 43.61 43.96 43.46 ;
      RECT  43.45 44.73 46.05 44.32 ;
      RECT  43.45 39.68 46.05 39.23 ;
      RECT  44.31 44.09 44.63 43.77 ;
      RECT  44.79 40.95 45.08 40.66 ;
      RECT  43.65 43.46 43.94 43.3 ;
      RECT  44.37 47.57 44.66 47.86 ;
      RECT  44.82 44.97 45.14 45.29 ;
      RECT  43.63 45.45 43.96 45.6 ;
      RECT  43.45 44.33 46.05 44.74 ;
      RECT  43.45 49.38 46.05 49.83 ;
      RECT  44.31 44.97 44.63 45.29 ;
      RECT  44.79 48.11 45.08 48.4 ;
      RECT  43.65 45.6 43.94 45.76 ;
      RECT  44.37 51.67 44.66 51.38 ;
      RECT  44.82 54.27 45.14 53.95 ;
      RECT  43.63 53.79 43.96 53.64 ;
      RECT  43.45 54.91 46.05 54.5 ;
      RECT  43.45 49.86 46.05 49.41 ;
      RECT  44.31 54.27 44.63 53.95 ;
      RECT  44.79 51.13 45.08 50.84 ;
      RECT  43.65 53.64 43.94 53.48 ;
      RECT  44.37 57.75 44.66 58.04 ;
      RECT  44.82 55.15 45.14 55.47 ;
      RECT  43.63 55.63 43.96 55.78 ;
      RECT  43.45 54.51 46.05 54.92 ;
      RECT  43.45 59.56 46.05 60.01 ;
      RECT  44.31 55.15 44.63 55.47 ;
      RECT  44.79 58.29 45.08 58.58 ;
      RECT  43.65 55.78 43.94 55.94 ;
      RECT  44.37 61.85 44.66 61.56 ;
      RECT  44.82 64.45 45.14 64.13 ;
      RECT  43.63 63.97 43.96 63.82 ;
      RECT  43.45 65.09 46.05 64.68 ;
      RECT  43.45 60.04 46.05 59.59 ;
      RECT  44.31 64.45 44.63 64.13 ;
      RECT  44.79 61.31 45.08 61.02 ;
      RECT  43.65 63.82 43.94 63.66 ;
      RECT  44.37 67.93 44.66 68.22 ;
      RECT  44.82 65.33 45.14 65.65 ;
      RECT  43.63 65.81 43.96 65.96 ;
      RECT  43.45 64.69 46.05 65.1 ;
      RECT  43.45 69.74 46.05 70.19 ;
      RECT  44.31 65.33 44.63 65.65 ;
      RECT  44.79 68.47 45.08 68.76 ;
      RECT  43.65 65.96 43.94 66.12 ;
      RECT  44.37 72.03 44.66 71.74 ;
      RECT  44.82 74.63 45.14 74.31 ;
      RECT  43.63 74.15 43.96 74.0 ;
      RECT  43.45 75.27 46.05 74.86 ;
      RECT  43.45 70.22 46.05 69.77 ;
      RECT  44.31 74.63 44.63 74.31 ;
      RECT  44.79 71.49 45.08 71.2 ;
      RECT  43.65 74.0 43.94 73.84 ;
      RECT  44.37 78.11 44.66 78.4 ;
      RECT  44.82 75.51 45.14 75.83 ;
      RECT  43.63 75.99 43.96 76.14 ;
      RECT  43.45 74.87 46.05 75.28 ;
      RECT  43.45 79.92 46.05 80.37 ;
      RECT  44.31 75.51 44.63 75.83 ;
      RECT  44.79 78.65 45.08 78.94 ;
      RECT  43.65 76.14 43.94 76.3 ;
      RECT  44.37 82.21 44.66 81.92 ;
      RECT  44.82 84.81 45.14 84.49 ;
      RECT  43.63 84.33 43.96 84.18 ;
      RECT  43.45 85.45 46.05 85.04 ;
      RECT  43.45 80.4 46.05 79.95 ;
      RECT  44.31 84.81 44.63 84.49 ;
      RECT  44.79 81.67 45.08 81.38 ;
      RECT  43.65 84.18 43.94 84.02 ;
      RECT  44.37 88.29 44.66 88.58 ;
      RECT  44.82 85.69 45.14 86.01 ;
      RECT  43.63 86.17 43.96 86.32 ;
      RECT  43.45 85.05 46.05 85.46 ;
      RECT  43.45 90.1 46.05 90.55 ;
      RECT  44.31 85.69 44.63 86.01 ;
      RECT  44.79 88.83 45.08 89.12 ;
      RECT  43.65 86.32 43.94 86.48 ;
      RECT  44.37 92.39 44.66 92.1 ;
      RECT  44.82 94.99 45.14 94.67 ;
      RECT  43.63 94.51 43.96 94.36 ;
      RECT  43.45 95.63 46.05 95.22 ;
      RECT  43.45 90.58 46.05 90.13 ;
      RECT  44.31 94.99 44.63 94.67 ;
      RECT  44.79 91.85 45.08 91.56 ;
      RECT  43.65 94.36 43.94 94.2 ;
      RECT  44.37 98.47 44.66 98.76 ;
      RECT  44.82 95.87 45.14 96.19 ;
      RECT  43.63 96.35 43.96 96.5 ;
      RECT  43.45 95.23 46.05 95.64 ;
      RECT  43.45 100.28 46.05 100.73 ;
      RECT  44.31 95.87 44.63 96.19 ;
      RECT  44.79 99.01 45.08 99.3 ;
      RECT  43.65 96.5 43.94 96.66 ;
      RECT  44.37 102.57 44.66 102.28 ;
      RECT  44.82 105.17 45.14 104.85 ;
      RECT  43.63 104.69 43.96 104.54 ;
      RECT  43.45 105.81 46.05 105.4 ;
      RECT  43.45 100.76 46.05 100.31 ;
      RECT  44.31 105.17 44.63 104.85 ;
      RECT  44.79 102.03 45.08 101.74 ;
      RECT  43.65 104.54 43.94 104.38 ;
      RECT  44.37 108.65 44.66 108.94 ;
      RECT  44.82 106.05 45.14 106.37 ;
      RECT  43.63 106.53 43.96 106.68 ;
      RECT  43.45 105.41 46.05 105.82 ;
      RECT  43.45 110.46 46.05 110.91 ;
      RECT  44.31 106.05 44.63 106.37 ;
      RECT  44.79 109.19 45.08 109.48 ;
      RECT  43.65 106.68 43.94 106.84 ;
      RECT  44.37 112.75 44.66 112.46 ;
      RECT  44.82 115.35 45.14 115.03 ;
      RECT  43.63 114.87 43.96 114.72 ;
      RECT  43.45 115.99 46.05 115.58 ;
      RECT  43.45 110.94 46.05 110.49 ;
      RECT  44.31 115.35 44.63 115.03 ;
      RECT  44.79 112.21 45.08 111.92 ;
      RECT  43.65 114.72 43.94 114.56 ;
      RECT  44.37 118.83 44.66 119.12 ;
      RECT  44.82 116.23 45.14 116.55 ;
      RECT  43.63 116.71 43.96 116.86 ;
      RECT  43.45 115.59 46.05 116.0 ;
      RECT  43.45 120.64 46.05 121.09 ;
      RECT  44.31 116.23 44.63 116.55 ;
      RECT  44.79 119.37 45.08 119.66 ;
      RECT  43.65 116.86 43.94 117.02 ;
      RECT  43.45 25.24 46.05 25.4 ;
      RECT  43.45 33.12 46.05 33.28 ;
      RECT  43.45 35.42 46.05 35.58 ;
      RECT  43.45 43.3 46.05 43.46 ;
      RECT  43.45 45.6 46.05 45.76 ;
      RECT  43.45 53.48 46.05 53.64 ;
      RECT  43.45 55.78 46.05 55.94 ;
      RECT  43.45 63.66 46.05 63.82 ;
      RECT  43.45 65.96 46.05 66.12 ;
      RECT  43.45 73.84 46.05 74.0 ;
      RECT  43.45 76.14 46.05 76.3 ;
      RECT  43.45 84.02 46.05 84.18 ;
      RECT  43.45 86.32 46.05 86.48 ;
      RECT  43.45 94.2 46.05 94.36 ;
      RECT  43.45 96.5 46.05 96.66 ;
      RECT  43.45 104.38 46.05 104.54 ;
      RECT  43.45 106.68 46.05 106.84 ;
      RECT  43.45 114.56 46.05 114.72 ;
      RECT  43.45 116.86 46.05 117.02 ;
      RECT  43.45 90.13 46.05 90.58 ;
      RECT  43.45 69.77 46.05 70.22 ;
      RECT  43.45 39.2 46.05 39.65 ;
      RECT  43.45 59.56 46.05 60.01 ;
      RECT  43.45 100.28 46.05 100.73 ;
      RECT  43.45 110.49 46.05 110.94 ;
      RECT  43.45 69.74 46.05 70.19 ;
      RECT  43.45 59.59 46.05 60.04 ;
      RECT  43.45 29.02 46.05 29.47 ;
      RECT  43.45 100.31 46.05 100.76 ;
      RECT  43.45 120.64 46.05 121.09 ;
      RECT  43.45 79.95 46.05 80.4 ;
      RECT  43.45 110.46 46.05 110.91 ;
      RECT  43.45 39.23 46.05 39.68 ;
      RECT  43.45 29.05 46.05 29.5 ;
      RECT  43.45 79.92 46.05 80.37 ;
      RECT  43.45 49.38 46.05 49.83 ;
      RECT  43.45 49.41 46.05 49.86 ;
      RECT  43.45 90.1 46.05 90.55 ;
      RECT  43.45 105.41 46.05 105.82 ;
      RECT  43.45 95.22 46.05 95.63 ;
      RECT  43.45 34.14 46.05 34.55 ;
      RECT  43.45 44.32 46.05 44.73 ;
      RECT  43.45 64.69 46.05 65.1 ;
      RECT  43.45 64.68 46.05 65.09 ;
      RECT  43.45 95.23 46.05 95.64 ;
      RECT  43.45 74.87 46.05 75.28 ;
      RECT  43.45 85.05 46.05 85.46 ;
      RECT  43.45 105.4 46.05 105.81 ;
      RECT  43.45 34.15 46.05 34.56 ;
      RECT  43.45 54.5 46.05 54.91 ;
      RECT  43.45 54.51 46.05 54.92 ;
      RECT  43.45 115.59 46.05 116.0 ;
      RECT  43.45 23.97 46.05 24.38 ;
      RECT  43.45 115.58 46.05 115.99 ;
      RECT  43.45 74.86 46.05 75.27 ;
      RECT  43.45 85.04 46.05 85.45 ;
      RECT  43.45 44.33 46.05 44.74 ;
      RECT  54.77 27.21 55.06 27.5 ;
      RECT  55.22 24.61 55.54 24.93 ;
      RECT  54.03 25.09 54.36 25.24 ;
      RECT  53.85 23.97 56.45 24.38 ;
      RECT  53.85 29.02 56.45 29.47 ;
      RECT  54.71 24.61 55.03 24.93 ;
      RECT  55.19 27.75 55.48 28.04 ;
      RECT  54.05 25.24 54.34 25.4 ;
      RECT  54.77 31.31 55.06 31.02 ;
      RECT  55.22 33.91 55.54 33.59 ;
      RECT  54.03 33.43 54.36 33.28 ;
      RECT  53.85 34.55 56.45 34.14 ;
      RECT  53.85 29.5 56.45 29.05 ;
      RECT  54.71 33.91 55.03 33.59 ;
      RECT  55.19 30.77 55.48 30.48 ;
      RECT  54.05 33.28 54.34 33.12 ;
      RECT  54.77 37.39 55.06 37.68 ;
      RECT  55.22 34.79 55.54 35.11 ;
      RECT  54.03 35.27 54.36 35.42 ;
      RECT  53.85 34.15 56.45 34.56 ;
      RECT  53.85 39.2 56.45 39.65 ;
      RECT  54.71 34.79 55.03 35.11 ;
      RECT  55.19 37.93 55.48 38.22 ;
      RECT  54.05 35.42 54.34 35.58 ;
      RECT  54.77 41.49 55.06 41.2 ;
      RECT  55.22 44.09 55.54 43.77 ;
      RECT  54.03 43.61 54.36 43.46 ;
      RECT  53.85 44.73 56.45 44.32 ;
      RECT  53.85 39.68 56.45 39.23 ;
      RECT  54.71 44.09 55.03 43.77 ;
      RECT  55.19 40.95 55.48 40.66 ;
      RECT  54.05 43.46 54.34 43.3 ;
      RECT  54.77 47.57 55.06 47.86 ;
      RECT  55.22 44.97 55.54 45.29 ;
      RECT  54.03 45.45 54.36 45.6 ;
      RECT  53.85 44.33 56.45 44.74 ;
      RECT  53.85 49.38 56.45 49.83 ;
      RECT  54.71 44.97 55.03 45.29 ;
      RECT  55.19 48.11 55.48 48.4 ;
      RECT  54.05 45.6 54.34 45.76 ;
      RECT  54.77 51.67 55.06 51.38 ;
      RECT  55.22 54.27 55.54 53.95 ;
      RECT  54.03 53.79 54.36 53.64 ;
      RECT  53.85 54.91 56.45 54.5 ;
      RECT  53.85 49.86 56.45 49.41 ;
      RECT  54.71 54.27 55.03 53.95 ;
      RECT  55.19 51.13 55.48 50.84 ;
      RECT  54.05 53.64 54.34 53.48 ;
      RECT  54.77 57.75 55.06 58.04 ;
      RECT  55.22 55.15 55.54 55.47 ;
      RECT  54.03 55.63 54.36 55.78 ;
      RECT  53.85 54.51 56.45 54.92 ;
      RECT  53.85 59.56 56.45 60.01 ;
      RECT  54.71 55.15 55.03 55.47 ;
      RECT  55.19 58.29 55.48 58.58 ;
      RECT  54.05 55.78 54.34 55.94 ;
      RECT  54.77 61.85 55.06 61.56 ;
      RECT  55.22 64.45 55.54 64.13 ;
      RECT  54.03 63.97 54.36 63.82 ;
      RECT  53.85 65.09 56.45 64.68 ;
      RECT  53.85 60.04 56.45 59.59 ;
      RECT  54.71 64.45 55.03 64.13 ;
      RECT  55.19 61.31 55.48 61.02 ;
      RECT  54.05 63.82 54.34 63.66 ;
      RECT  54.77 67.93 55.06 68.22 ;
      RECT  55.22 65.33 55.54 65.65 ;
      RECT  54.03 65.81 54.36 65.96 ;
      RECT  53.85 64.69 56.45 65.1 ;
      RECT  53.85 69.74 56.45 70.19 ;
      RECT  54.71 65.33 55.03 65.65 ;
      RECT  55.19 68.47 55.48 68.76 ;
      RECT  54.05 65.96 54.34 66.12 ;
      RECT  54.77 72.03 55.06 71.74 ;
      RECT  55.22 74.63 55.54 74.31 ;
      RECT  54.03 74.15 54.36 74.0 ;
      RECT  53.85 75.27 56.45 74.86 ;
      RECT  53.85 70.22 56.45 69.77 ;
      RECT  54.71 74.63 55.03 74.31 ;
      RECT  55.19 71.49 55.48 71.2 ;
      RECT  54.05 74.0 54.34 73.84 ;
      RECT  54.77 78.11 55.06 78.4 ;
      RECT  55.22 75.51 55.54 75.83 ;
      RECT  54.03 75.99 54.36 76.14 ;
      RECT  53.85 74.87 56.45 75.28 ;
      RECT  53.85 79.92 56.45 80.37 ;
      RECT  54.71 75.51 55.03 75.83 ;
      RECT  55.19 78.65 55.48 78.94 ;
      RECT  54.05 76.14 54.34 76.3 ;
      RECT  54.77 82.21 55.06 81.92 ;
      RECT  55.22 84.81 55.54 84.49 ;
      RECT  54.03 84.33 54.36 84.18 ;
      RECT  53.85 85.45 56.45 85.04 ;
      RECT  53.85 80.4 56.45 79.95 ;
      RECT  54.71 84.81 55.03 84.49 ;
      RECT  55.19 81.67 55.48 81.38 ;
      RECT  54.05 84.18 54.34 84.02 ;
      RECT  54.77 88.29 55.06 88.58 ;
      RECT  55.22 85.69 55.54 86.01 ;
      RECT  54.03 86.17 54.36 86.32 ;
      RECT  53.85 85.05 56.45 85.46 ;
      RECT  53.85 90.1 56.45 90.55 ;
      RECT  54.71 85.69 55.03 86.01 ;
      RECT  55.19 88.83 55.48 89.12 ;
      RECT  54.05 86.32 54.34 86.48 ;
      RECT  54.77 92.39 55.06 92.1 ;
      RECT  55.22 94.99 55.54 94.67 ;
      RECT  54.03 94.51 54.36 94.36 ;
      RECT  53.85 95.63 56.45 95.22 ;
      RECT  53.85 90.58 56.45 90.13 ;
      RECT  54.71 94.99 55.03 94.67 ;
      RECT  55.19 91.85 55.48 91.56 ;
      RECT  54.05 94.36 54.34 94.2 ;
      RECT  54.77 98.47 55.06 98.76 ;
      RECT  55.22 95.87 55.54 96.19 ;
      RECT  54.03 96.35 54.36 96.5 ;
      RECT  53.85 95.23 56.45 95.64 ;
      RECT  53.85 100.28 56.45 100.73 ;
      RECT  54.71 95.87 55.03 96.19 ;
      RECT  55.19 99.01 55.48 99.3 ;
      RECT  54.05 96.5 54.34 96.66 ;
      RECT  54.77 102.57 55.06 102.28 ;
      RECT  55.22 105.17 55.54 104.85 ;
      RECT  54.03 104.69 54.36 104.54 ;
      RECT  53.85 105.81 56.45 105.4 ;
      RECT  53.85 100.76 56.45 100.31 ;
      RECT  54.71 105.17 55.03 104.85 ;
      RECT  55.19 102.03 55.48 101.74 ;
      RECT  54.05 104.54 54.34 104.38 ;
      RECT  54.77 108.65 55.06 108.94 ;
      RECT  55.22 106.05 55.54 106.37 ;
      RECT  54.03 106.53 54.36 106.68 ;
      RECT  53.85 105.41 56.45 105.82 ;
      RECT  53.85 110.46 56.45 110.91 ;
      RECT  54.71 106.05 55.03 106.37 ;
      RECT  55.19 109.19 55.48 109.48 ;
      RECT  54.05 106.68 54.34 106.84 ;
      RECT  54.77 112.75 55.06 112.46 ;
      RECT  55.22 115.35 55.54 115.03 ;
      RECT  54.03 114.87 54.36 114.72 ;
      RECT  53.85 115.99 56.45 115.58 ;
      RECT  53.85 110.94 56.45 110.49 ;
      RECT  54.71 115.35 55.03 115.03 ;
      RECT  55.19 112.21 55.48 111.92 ;
      RECT  54.05 114.72 54.34 114.56 ;
      RECT  54.77 118.83 55.06 119.12 ;
      RECT  55.22 116.23 55.54 116.55 ;
      RECT  54.03 116.71 54.36 116.86 ;
      RECT  53.85 115.59 56.45 116.0 ;
      RECT  53.85 120.64 56.45 121.09 ;
      RECT  54.71 116.23 55.03 116.55 ;
      RECT  55.19 119.37 55.48 119.66 ;
      RECT  54.05 116.86 54.34 117.02 ;
      RECT  53.85 25.24 56.45 25.4 ;
      RECT  53.85 33.12 56.45 33.28 ;
      RECT  53.85 35.42 56.45 35.58 ;
      RECT  53.85 43.3 56.45 43.46 ;
      RECT  53.85 45.6 56.45 45.76 ;
      RECT  53.85 53.48 56.45 53.64 ;
      RECT  53.85 55.78 56.45 55.94 ;
      RECT  53.85 63.66 56.45 63.82 ;
      RECT  53.85 65.96 56.45 66.12 ;
      RECT  53.85 73.84 56.45 74.0 ;
      RECT  53.85 76.14 56.45 76.3 ;
      RECT  53.85 84.02 56.45 84.18 ;
      RECT  53.85 86.32 56.45 86.48 ;
      RECT  53.85 94.2 56.45 94.36 ;
      RECT  53.85 96.5 56.45 96.66 ;
      RECT  53.85 104.38 56.45 104.54 ;
      RECT  53.85 106.68 56.45 106.84 ;
      RECT  53.85 114.56 56.45 114.72 ;
      RECT  53.85 116.86 56.45 117.02 ;
      RECT  53.85 90.13 56.45 90.58 ;
      RECT  53.85 69.77 56.45 70.22 ;
      RECT  53.85 39.2 56.45 39.65 ;
      RECT  53.85 59.56 56.45 60.01 ;
      RECT  53.85 100.28 56.45 100.73 ;
      RECT  53.85 110.49 56.45 110.94 ;
      RECT  53.85 69.74 56.45 70.19 ;
      RECT  53.85 59.59 56.45 60.04 ;
      RECT  53.85 29.02 56.45 29.47 ;
      RECT  53.85 100.31 56.45 100.76 ;
      RECT  53.85 120.64 56.45 121.09 ;
      RECT  53.85 79.95 56.45 80.4 ;
      RECT  53.85 110.46 56.45 110.91 ;
      RECT  53.85 39.23 56.45 39.68 ;
      RECT  53.85 29.05 56.45 29.5 ;
      RECT  53.85 79.92 56.45 80.37 ;
      RECT  53.85 49.38 56.45 49.83 ;
      RECT  53.85 49.41 56.45 49.86 ;
      RECT  53.85 90.1 56.45 90.55 ;
      RECT  53.85 105.41 56.45 105.82 ;
      RECT  53.85 95.22 56.45 95.63 ;
      RECT  53.85 34.14 56.45 34.55 ;
      RECT  53.85 44.32 56.45 44.73 ;
      RECT  53.85 64.69 56.45 65.1 ;
      RECT  53.85 64.68 56.45 65.09 ;
      RECT  53.85 95.23 56.45 95.64 ;
      RECT  53.85 74.87 56.45 75.28 ;
      RECT  53.85 85.05 56.45 85.46 ;
      RECT  53.85 105.4 56.45 105.81 ;
      RECT  53.85 34.15 56.45 34.56 ;
      RECT  53.85 54.5 56.45 54.91 ;
      RECT  53.85 54.51 56.45 54.92 ;
      RECT  53.85 115.59 56.45 116.0 ;
      RECT  53.85 23.97 56.45 24.38 ;
      RECT  53.85 115.58 56.45 115.99 ;
      RECT  53.85 74.86 56.45 75.27 ;
      RECT  53.85 85.04 56.45 85.45 ;
      RECT  53.85 44.33 56.45 44.74 ;
      RECT  42.55 33.12 57.35 33.28 ;
      RECT  42.55 35.42 57.35 35.58 ;
      RECT  42.55 43.3 57.35 43.46 ;
      RECT  42.55 45.6 57.35 45.76 ;
      RECT  42.55 53.48 57.35 53.64 ;
      RECT  42.55 55.78 57.35 55.94 ;
      RECT  42.55 63.66 57.35 63.82 ;
      RECT  42.55 65.96 57.35 66.12 ;
      RECT  42.55 73.84 57.35 74.0 ;
      RECT  42.55 76.14 57.35 76.3 ;
      RECT  42.55 84.02 57.35 84.18 ;
      RECT  42.55 86.32 57.35 86.48 ;
      RECT  42.55 94.2 57.35 94.36 ;
      RECT  42.55 96.5 57.35 96.66 ;
      RECT  42.55 104.38 57.35 104.54 ;
      RECT  42.55 106.68 57.35 106.84 ;
      RECT  42.55 114.56 57.35 114.72 ;
      RECT  46.05 90.13 48.65 90.58 ;
      RECT  46.05 59.56 48.65 60.01 ;
      RECT  46.05 59.59 48.65 60.04 ;
      RECT  46.05 110.46 48.65 110.91 ;
      RECT  46.05 79.95 48.65 80.4 ;
      RECT  46.05 90.1 48.65 90.55 ;
      RECT  46.05 100.28 48.65 100.73 ;
      RECT  46.05 79.92 48.65 80.37 ;
      RECT  46.05 69.77 48.65 70.22 ;
      RECT  46.05 110.49 48.65 110.94 ;
      RECT  46.05 49.41 48.65 49.86 ;
      RECT  46.05 39.23 48.65 39.68 ;
      RECT  46.05 39.2 48.65 39.65 ;
      RECT  46.05 49.38 48.65 49.83 ;
      RECT  46.05 100.31 48.65 100.76 ;
      RECT  46.05 69.74 48.65 70.19 ;
      RECT  46.05 29.05 48.65 29.5 ;
      RECT  46.05 64.68 48.65 65.09 ;
      RECT  46.05 74.86 48.65 75.27 ;
      RECT  46.05 54.5 48.65 54.91 ;
      RECT  46.05 74.87 48.65 75.28 ;
      RECT  46.05 95.23 48.65 95.64 ;
      RECT  46.05 44.33 48.65 44.74 ;
      RECT  46.05 105.41 48.65 105.82 ;
      RECT  46.05 95.22 48.65 95.63 ;
      RECT  46.05 105.4 48.65 105.81 ;
      RECT  46.05 34.14 48.65 34.55 ;
      RECT  46.05 64.69 48.65 65.1 ;
      RECT  46.05 44.32 48.65 44.73 ;
      RECT  46.05 115.58 48.65 115.99 ;
      RECT  46.05 85.05 48.65 85.46 ;
      RECT  46.05 54.51 48.65 54.92 ;
      RECT  46.05 85.04 48.65 85.45 ;
      RECT  46.05 34.15 48.65 34.56 ;
      RECT  46.05 16.35 48.65 16.49 ;
      RECT  48.65 16.35 51.25 16.49 ;
      RECT  51.25 16.35 53.85 16.49 ;
      RECT  42.55 16.35 53.85 16.49 ;
      RECT  48.82 10.6 52.09 10.89 ;
      RECT  53.94 10.57 54.27 11.17 ;
      RECT  50.0 9.64 50.33 10.28 ;
      RECT  48.35 8.63 54.42 9.04 ;
      RECT  53.09 9.9 54.42 10.23 ;
      RECT  48.35 9.62 48.69 10.28 ;
      RECT  48.35 13.0 54.42 13.41 ;
      RECT  51.42 10.6 54.69 10.89 ;
      RECT  56.54 10.57 56.87 11.17 ;
      RECT  52.6 9.64 52.93 10.28 ;
      RECT  50.95 8.63 57.02 9.04 ;
      RECT  55.69 9.9 57.02 10.23 ;
      RECT  50.95 9.62 51.29 10.28 ;
      RECT  50.95 13.0 57.02 13.41 ;
      RECT  42.55 9.99 57.02 10.13 ;
      RECT  51.42 3.55 51.72 3.6 ;
      RECT  49.82 6.94 62.06 7.39 ;
      RECT  51.42 3.8 51.72 3.85 ;
      RECT  59.59 3.97 59.92 4.01 ;
      RECT  53.73 3.08 54.03 5.7 ;
      RECT  60.04 5.41 60.34 5.7 ;
      RECT  49.82 1.15 62.06 1.57 ;
      RECT  60.08 3.37 60.34 5.41 ;
      RECT  60.04 3.08 60.34 3.37 ;
      RECT  61.59 4.41 61.89 4.7 ;
      RECT  61.75 3.04 62.05 3.33 ;
      RECT  49.82 3.6 51.72 3.8 ;
      RECT  49.92 3.02 50.25 3.35 ;
      RECT  54.98 3.68 59.92 3.97 ;
      RECT  55.43 4.41 59.26 4.7 ;
      RECT  54.02 3.55 54.32 3.6 ;
      RECT  52.42 6.94 64.66 7.39 ;
      RECT  54.02 3.8 54.32 3.85 ;
      RECT  62.19 3.97 62.52 4.01 ;
      RECT  56.33 3.08 56.63 5.7 ;
      RECT  62.64 5.41 62.94 5.7 ;
      RECT  52.42 1.15 64.66 1.57 ;
      RECT  62.68 3.37 62.94 5.41 ;
      RECT  62.64 3.08 62.94 3.37 ;
      RECT  64.19 4.41 64.49 4.7 ;
      RECT  64.35 3.04 64.65 3.33 ;
      RECT  52.42 3.6 54.32 3.8 ;
      RECT  52.52 3.02 52.85 3.35 ;
      RECT  57.58 3.68 62.52 3.97 ;
      RECT  58.03 4.41 61.86 4.7 ;
      RECT  42.55 3.68 64.66 3.82 ;
      RECT  42.55 10.13 57.02 9.99 ;
      RECT  42.55 16.49 53.85 16.35 ;
      RECT  42.55 3.82 64.66 3.68 ;
      RECT  -53.04 -7.17 -52.71 -7.16 ;
      RECT  -55.28 -8.11 -53.83 -7.91 ;
      RECT  -53.04 -7.41 -52.71 -7.38 ;
      RECT  -47.24 -7.17 -46.91 -7.16 ;
      RECT  -56.23 -5.67 -43.52 -5.22 ;
      RECT  -55.28 -7.91 -54.99 -7.85 ;
      RECT  -46.1 -7.51 -45.47 -7.19 ;
      RECT  -48.32 -7.83 -48.12 -7.66 ;
      RECT  -48.32 -7.41 -48.12 -7.16 ;
      RECT  -47.63 -8.26 -44.1 -8.06 ;
      RECT  -53.04 -7.66 -48.12 -7.41 ;
      RECT  -54.12 -7.16 -48.63 -6.96 ;
      RECT  -54.16 -8.16 -53.83 -8.11 ;
      RECT  -56.15 -8.02 -55.47 -7.7 ;
      RECT  -48.96 -7.17 -48.63 -7.16 ;
      RECT  -54.16 -7.91 -53.83 -7.83 ;
      RECT  -56.23 -9.76 -43.52 -9.31 ;
      RECT  -44.44 -8.36 -44.1 -8.26 ;
      RECT  -53.04 -6.96 -52.71 -6.84 ;
      RECT  -44.44 -8.06 -44.1 -8.03 ;
      RECT  -54.12 -7.83 -53.92 -7.16 ;
      RECT  -48.32 -7.16 -46.91 -6.96 ;
      RECT  -48.96 -6.96 -48.63 -6.84 ;
      RECT  -48.36 -8.16 -48.03 -7.83 ;
      RECT  -53.43 -8.06 -53.13 -7.96 ;
      RECT  -50.47 -8.32 -50.14 -8.27 ;
      RECT  -55.0 -7.2 -54.37 -6.88 ;
      RECT  -53.43 -8.27 -50.14 -8.06 ;
      RECT  -47.63 -8.06 -47.33 -7.95 ;
      RECT  -47.24 -6.96 -46.91 -6.84 ;
      RECT  -53.04 -7.71 -52.71 -7.66 ;
      RECT  -50.47 -8.06 -50.14 -7.99 ;
      RECT  -55.28 -8.14 -54.99 -8.11 ;
      RECT  -56.23 -5.67 -33.42 -5.22 ;
      RECT  -56.23 -9.76 -33.42 -9.31 ;
      RECT  -53.04 -3.73 -52.71 -3.74 ;
      RECT  -55.28 -2.79 -53.83 -2.99 ;
      RECT  -53.04 -3.49 -52.71 -3.52 ;
      RECT  -47.24 -3.73 -46.91 -3.74 ;
      RECT  -56.23 -5.23 -43.52 -5.68 ;
      RECT  -55.28 -2.99 -54.99 -3.05 ;
      RECT  -46.1 -3.39 -45.47 -3.71 ;
      RECT  -48.32 -3.07 -48.12 -3.24 ;
      RECT  -48.32 -3.49 -48.12 -3.74 ;
      RECT  -47.63 -2.64 -44.1 -2.84 ;
      RECT  -53.04 -3.24 -48.12 -3.49 ;
      RECT  -54.12 -3.74 -48.63 -3.94 ;
      RECT  -54.16 -2.74 -53.83 -2.79 ;
      RECT  -56.15 -2.88 -55.47 -3.2 ;
      RECT  -48.96 -3.73 -48.63 -3.74 ;
      RECT  -54.16 -2.99 -53.83 -3.07 ;
      RECT  -56.23 -1.14 -43.52 -1.59 ;
      RECT  -44.44 -2.54 -44.1 -2.64 ;
      RECT  -53.04 -3.94 -52.71 -4.06 ;
      RECT  -44.44 -2.84 -44.1 -2.87 ;
      RECT  -54.12 -3.07 -53.92 -3.74 ;
      RECT  -48.32 -3.74 -46.91 -3.94 ;
      RECT  -48.96 -3.94 -48.63 -4.06 ;
      RECT  -48.36 -2.74 -48.03 -3.07 ;
      RECT  -53.43 -2.84 -53.13 -2.94 ;
      RECT  -50.47 -2.58 -50.14 -2.63 ;
      RECT  -55.0 -3.7 -54.37 -4.02 ;
      RECT  -53.43 -2.63 -50.14 -2.84 ;
      RECT  -47.63 -2.84 -47.33 -2.95 ;
      RECT  -47.24 -3.94 -46.91 -4.06 ;
      RECT  -53.04 -3.19 -52.71 -3.24 ;
      RECT  -50.47 -2.84 -50.14 -2.91 ;
      RECT  -55.28 -2.76 -54.99 -2.79 ;
      RECT  -56.23 -5.23 -33.42 -5.68 ;
      RECT  -56.23 -1.14 -33.42 -1.59 ;
      RECT  -10.84 103.31 -10.51 103.32 ;
      RECT  -13.08 102.37 -11.63 102.57 ;
      RECT  -10.84 103.07 -10.51 103.1 ;
      RECT  -5.04 103.31 -4.71 103.32 ;
      RECT  -14.03 104.81 -1.32 105.26 ;
      RECT  -13.08 102.57 -12.79 102.63 ;
      RECT  -3.9 102.97 -3.27 103.29 ;
      RECT  -6.12 102.65 -5.92 102.82 ;
      RECT  -6.12 103.07 -5.92 103.32 ;
      RECT  -5.43 102.22 -1.9 102.42 ;
      RECT  -10.84 102.82 -5.92 103.07 ;
      RECT  -11.92 103.32 -6.43 103.52 ;
      RECT  -11.96 102.32 -11.63 102.37 ;
      RECT  -13.95 102.46 -13.27 102.78 ;
      RECT  -6.76 103.31 -6.43 103.32 ;
      RECT  -11.96 102.57 -11.63 102.65 ;
      RECT  -14.03 100.72 -1.32 101.17 ;
      RECT  -2.24 102.12 -1.9 102.22 ;
      RECT  -10.84 103.52 -10.51 103.64 ;
      RECT  -2.24 102.42 -1.9 102.45 ;
      RECT  -11.92 102.65 -11.72 103.32 ;
      RECT  -6.12 103.32 -4.71 103.52 ;
      RECT  -6.76 103.52 -6.43 103.64 ;
      RECT  -6.16 102.32 -5.83 102.65 ;
      RECT  -11.23 102.42 -10.93 102.52 ;
      RECT  -8.27 102.16 -7.94 102.21 ;
      RECT  -12.8 103.28 -12.17 103.6 ;
      RECT  -11.23 102.21 -7.94 102.42 ;
      RECT  -5.43 102.42 -5.13 102.53 ;
      RECT  -5.04 103.52 -4.71 103.64 ;
      RECT  -10.84 102.77 -10.51 102.82 ;
      RECT  -8.27 102.42 -7.94 102.49 ;
      RECT  -13.08 102.34 -12.79 102.37 ;
      RECT  -10.84 106.75 -10.51 106.74 ;
      RECT  -13.08 107.69 -11.63 107.49 ;
      RECT  -10.84 106.99 -10.51 106.96 ;
      RECT  -5.04 106.75 -4.71 106.74 ;
      RECT  -14.03 105.25 -1.32 104.8 ;
      RECT  -13.08 107.49 -12.79 107.43 ;
      RECT  -3.9 107.09 -3.27 106.77 ;
      RECT  -6.12 107.41 -5.92 107.24 ;
      RECT  -6.12 106.99 -5.92 106.74 ;
      RECT  -5.43 107.84 -1.9 107.64 ;
      RECT  -10.84 107.24 -5.92 106.99 ;
      RECT  -11.92 106.74 -6.43 106.54 ;
      RECT  -11.96 107.74 -11.63 107.69 ;
      RECT  -13.95 107.6 -13.27 107.28 ;
      RECT  -6.76 106.75 -6.43 106.74 ;
      RECT  -11.96 107.49 -11.63 107.41 ;
      RECT  -14.03 109.34 -1.32 108.89 ;
      RECT  -2.24 107.94 -1.9 107.84 ;
      RECT  -10.84 106.54 -10.51 106.42 ;
      RECT  -2.24 107.64 -1.9 107.61 ;
      RECT  -11.92 107.41 -11.72 106.74 ;
      RECT  -6.12 106.74 -4.71 106.54 ;
      RECT  -6.76 106.54 -6.43 106.42 ;
      RECT  -6.16 107.74 -5.83 107.41 ;
      RECT  -11.23 107.64 -10.93 107.54 ;
      RECT  -8.27 107.9 -7.94 107.85 ;
      RECT  -12.8 106.78 -12.17 106.46 ;
      RECT  -11.23 107.85 -7.94 107.64 ;
      RECT  -5.43 107.64 -5.13 107.53 ;
      RECT  -5.04 106.54 -4.71 106.42 ;
      RECT  -10.84 107.29 -10.51 107.24 ;
      RECT  -8.27 107.64 -7.94 107.57 ;
      RECT  -13.08 107.72 -12.79 107.69 ;
      RECT  -10.84 111.43 -10.51 111.44 ;
      RECT  -13.08 110.49 -11.63 110.69 ;
      RECT  -10.84 111.19 -10.51 111.22 ;
      RECT  -5.04 111.43 -4.71 111.44 ;
      RECT  -14.03 112.93 -1.32 113.38 ;
      RECT  -13.08 110.69 -12.79 110.75 ;
      RECT  -3.9 111.09 -3.27 111.41 ;
      RECT  -6.12 110.77 -5.92 110.94 ;
      RECT  -6.12 111.19 -5.92 111.44 ;
      RECT  -5.43 110.34 -1.9 110.54 ;
      RECT  -10.84 110.94 -5.92 111.19 ;
      RECT  -11.92 111.44 -6.43 111.64 ;
      RECT  -11.96 110.44 -11.63 110.49 ;
      RECT  -13.95 110.58 -13.27 110.9 ;
      RECT  -6.76 111.43 -6.43 111.44 ;
      RECT  -11.96 110.69 -11.63 110.77 ;
      RECT  -14.03 108.84 -1.32 109.29 ;
      RECT  -2.24 110.24 -1.9 110.34 ;
      RECT  -10.84 111.64 -10.51 111.76 ;
      RECT  -2.24 110.54 -1.9 110.57 ;
      RECT  -11.92 110.77 -11.72 111.44 ;
      RECT  -6.12 111.44 -4.71 111.64 ;
      RECT  -6.76 111.64 -6.43 111.76 ;
      RECT  -6.16 110.44 -5.83 110.77 ;
      RECT  -11.23 110.54 -10.93 110.64 ;
      RECT  -8.27 110.28 -7.94 110.33 ;
      RECT  -12.8 111.4 -12.17 111.72 ;
      RECT  -11.23 110.33 -7.94 110.54 ;
      RECT  -5.43 110.54 -5.13 110.65 ;
      RECT  -5.04 111.64 -4.71 111.76 ;
      RECT  -10.84 110.89 -10.51 110.94 ;
      RECT  -8.27 110.54 -7.94 110.61 ;
      RECT  -13.08 110.46 -12.79 110.49 ;
      RECT  -10.84 114.87 -10.51 114.86 ;
      RECT  -13.08 115.81 -11.63 115.61 ;
      RECT  -10.84 115.11 -10.51 115.08 ;
      RECT  -5.04 114.87 -4.71 114.86 ;
      RECT  -14.03 113.37 -1.32 112.92 ;
      RECT  -13.08 115.61 -12.79 115.55 ;
      RECT  -3.9 115.21 -3.27 114.89 ;
      RECT  -6.12 115.53 -5.92 115.36 ;
      RECT  -6.12 115.11 -5.92 114.86 ;
      RECT  -5.43 115.96 -1.9 115.76 ;
      RECT  -10.84 115.36 -5.92 115.11 ;
      RECT  -11.92 114.86 -6.43 114.66 ;
      RECT  -11.96 115.86 -11.63 115.81 ;
      RECT  -13.95 115.72 -13.27 115.4 ;
      RECT  -6.76 114.87 -6.43 114.86 ;
      RECT  -11.96 115.61 -11.63 115.53 ;
      RECT  -14.03 117.46 -1.32 117.01 ;
      RECT  -2.24 116.06 -1.9 115.96 ;
      RECT  -10.84 114.66 -10.51 114.54 ;
      RECT  -2.24 115.76 -1.9 115.73 ;
      RECT  -11.92 115.53 -11.72 114.86 ;
      RECT  -6.12 114.86 -4.71 114.66 ;
      RECT  -6.76 114.66 -6.43 114.54 ;
      RECT  -6.16 115.86 -5.83 115.53 ;
      RECT  -11.23 115.76 -10.93 115.66 ;
      RECT  -8.27 116.02 -7.94 115.97 ;
      RECT  -12.8 114.9 -12.17 114.58 ;
      RECT  -11.23 115.97 -7.94 115.76 ;
      RECT  -5.43 115.76 -5.13 115.65 ;
      RECT  -5.04 114.66 -4.71 114.54 ;
      RECT  -10.84 115.41 -10.51 115.36 ;
      RECT  -8.27 115.76 -7.94 115.69 ;
      RECT  -13.08 115.84 -12.79 115.81 ;
      RECT  12.46 -7.17 12.79 -7.16 ;
      RECT  10.22 -8.11 11.67 -7.91 ;
      RECT  12.46 -7.41 12.79 -7.38 ;
      RECT  18.26 -7.17 18.59 -7.16 ;
      RECT  9.27 -5.67 21.98 -5.22 ;
      RECT  10.22 -7.91 10.51 -7.85 ;
      RECT  19.4 -7.51 20.03 -7.19 ;
      RECT  17.18 -7.83 17.38 -7.66 ;
      RECT  17.18 -7.41 17.38 -7.16 ;
      RECT  17.87 -8.26 21.4 -8.06 ;
      RECT  12.46 -7.66 17.38 -7.41 ;
      RECT  11.38 -7.16 16.87 -6.96 ;
      RECT  11.34 -8.16 11.67 -8.11 ;
      RECT  9.35 -8.02 10.03 -7.7 ;
      RECT  16.54 -7.17 16.87 -7.16 ;
      RECT  11.34 -7.91 11.67 -7.83 ;
      RECT  9.27 -9.76 21.98 -9.31 ;
      RECT  21.06 -8.36 21.4 -8.26 ;
      RECT  12.46 -6.96 12.79 -6.84 ;
      RECT  21.06 -8.06 21.4 -8.03 ;
      RECT  11.38 -7.83 11.58 -7.16 ;
      RECT  17.18 -7.16 18.59 -6.96 ;
      RECT  16.54 -6.96 16.87 -6.84 ;
      RECT  17.14 -8.16 17.47 -7.83 ;
      RECT  12.07 -8.06 12.37 -7.96 ;
      RECT  15.03 -8.32 15.36 -8.27 ;
      RECT  10.5 -7.2 11.13 -6.88 ;
      RECT  12.07 -8.27 15.36 -8.06 ;
      RECT  17.87 -8.06 18.17 -7.95 ;
      RECT  18.26 -6.96 18.59 -6.84 ;
      RECT  12.46 -7.71 12.79 -7.66 ;
      RECT  15.03 -8.06 15.36 -7.99 ;
      RECT  10.22 -8.14 10.51 -8.11 ;
      RECT  24.11 -7.17 24.44 -7.16 ;
      RECT  21.87 -8.11 23.32 -7.91 ;
      RECT  24.11 -7.41 24.44 -7.38 ;
      RECT  29.91 -7.17 30.24 -7.16 ;
      RECT  20.92 -5.67 33.63 -5.22 ;
      RECT  21.87 -7.91 22.16 -7.85 ;
      RECT  31.05 -7.51 31.68 -7.19 ;
      RECT  28.83 -7.83 29.03 -7.66 ;
      RECT  28.83 -7.41 29.03 -7.16 ;
      RECT  29.52 -8.26 33.05 -8.06 ;
      RECT  24.11 -7.66 29.03 -7.41 ;
      RECT  23.03 -7.16 28.52 -6.96 ;
      RECT  22.99 -8.16 23.32 -8.11 ;
      RECT  21.0 -8.02 21.68 -7.7 ;
      RECT  28.19 -7.17 28.52 -7.16 ;
      RECT  22.99 -7.91 23.32 -7.83 ;
      RECT  20.92 -9.76 33.63 -9.31 ;
      RECT  32.71 -8.36 33.05 -8.26 ;
      RECT  24.11 -6.96 24.44 -6.84 ;
      RECT  32.71 -8.06 33.05 -8.03 ;
      RECT  23.03 -7.83 23.23 -7.16 ;
      RECT  28.83 -7.16 30.24 -6.96 ;
      RECT  28.19 -6.96 28.52 -6.84 ;
      RECT  28.79 -8.16 29.12 -7.83 ;
      RECT  23.72 -8.06 24.02 -7.96 ;
      RECT  26.68 -8.32 27.01 -8.27 ;
      RECT  22.15 -7.2 22.78 -6.88 ;
      RECT  23.72 -8.27 27.01 -8.06 ;
      RECT  29.52 -8.06 29.82 -7.95 ;
      RECT  29.91 -6.96 30.24 -6.84 ;
      RECT  24.11 -7.71 24.44 -7.66 ;
      RECT  26.68 -8.06 27.01 -7.99 ;
      RECT  21.87 -8.14 22.16 -8.11 ;
   LAYER  m2 ;
      RECT  50.02 34.87 50.74 35.01 ;
      RECT  49.51 34.79 49.83 34.86 ;
      RECT  49.51 35.0 49.83 35.11 ;
      RECT  50.02 35.01 50.34 35.11 ;
      RECT  49.18 35.0 49.32 39.89 ;
      RECT  50.6 34.15 50.74 34.87 ;
      RECT  49.18 34.15 49.32 34.86 ;
      RECT  50.6 35.01 50.74 39.89 ;
      RECT  50.02 34.79 50.34 34.87 ;
      RECT  49.18 34.86 49.83 35.0 ;
      RECT  50.02 44.01 50.74 43.87 ;
      RECT  49.51 44.09 49.83 44.02 ;
      RECT  49.51 43.88 49.83 43.77 ;
      RECT  50.02 43.87 50.34 43.77 ;
      RECT  49.18 43.88 49.32 38.99 ;
      RECT  50.6 44.73 50.74 44.01 ;
      RECT  49.18 44.73 49.32 44.02 ;
      RECT  50.6 43.87 50.74 38.99 ;
      RECT  50.02 44.09 50.34 44.01 ;
      RECT  49.18 44.02 49.83 43.88 ;
      RECT  50.02 45.05 50.74 45.19 ;
      RECT  49.51 44.97 49.83 45.04 ;
      RECT  49.51 45.18 49.83 45.29 ;
      RECT  50.02 45.19 50.34 45.29 ;
      RECT  49.18 45.18 49.32 50.07 ;
      RECT  50.6 44.33 50.74 45.05 ;
      RECT  49.18 44.33 49.32 45.04 ;
      RECT  50.6 45.19 50.74 50.07 ;
      RECT  50.02 44.97 50.34 45.05 ;
      RECT  49.18 45.04 49.83 45.18 ;
      RECT  50.02 54.19 50.74 54.05 ;
      RECT  49.51 54.27 49.83 54.2 ;
      RECT  49.51 54.06 49.83 53.95 ;
      RECT  50.02 54.05 50.34 53.95 ;
      RECT  49.18 54.06 49.32 49.17 ;
      RECT  50.6 54.91 50.74 54.19 ;
      RECT  49.18 54.91 49.32 54.2 ;
      RECT  50.6 54.05 50.74 49.17 ;
      RECT  50.02 54.27 50.34 54.19 ;
      RECT  49.18 54.2 49.83 54.06 ;
      RECT  50.02 55.23 50.74 55.37 ;
      RECT  49.51 55.15 49.83 55.22 ;
      RECT  49.51 55.36 49.83 55.47 ;
      RECT  50.02 55.37 50.34 55.47 ;
      RECT  49.18 55.36 49.32 60.25 ;
      RECT  50.6 54.51 50.74 55.23 ;
      RECT  49.18 54.51 49.32 55.22 ;
      RECT  50.6 55.37 50.74 60.25 ;
      RECT  50.02 55.15 50.34 55.23 ;
      RECT  49.18 55.22 49.83 55.36 ;
      RECT  50.02 64.37 50.74 64.23 ;
      RECT  49.51 64.45 49.83 64.38 ;
      RECT  49.51 64.24 49.83 64.13 ;
      RECT  50.02 64.23 50.34 64.13 ;
      RECT  49.18 64.24 49.32 59.35 ;
      RECT  50.6 65.09 50.74 64.37 ;
      RECT  49.18 65.09 49.32 64.38 ;
      RECT  50.6 64.23 50.74 59.35 ;
      RECT  50.02 64.45 50.34 64.37 ;
      RECT  49.18 64.38 49.83 64.24 ;
      RECT  50.02 65.41 50.74 65.55 ;
      RECT  49.51 65.33 49.83 65.4 ;
      RECT  49.51 65.54 49.83 65.65 ;
      RECT  50.02 65.55 50.34 65.65 ;
      RECT  49.18 65.54 49.32 70.43 ;
      RECT  50.6 64.69 50.74 65.41 ;
      RECT  49.18 64.69 49.32 65.4 ;
      RECT  50.6 65.55 50.74 70.43 ;
      RECT  50.02 65.33 50.34 65.41 ;
      RECT  49.18 65.4 49.83 65.54 ;
      RECT  50.02 74.55 50.74 74.41 ;
      RECT  49.51 74.63 49.83 74.56 ;
      RECT  49.51 74.42 49.83 74.31 ;
      RECT  50.02 74.41 50.34 74.31 ;
      RECT  49.18 74.42 49.32 69.53 ;
      RECT  50.6 75.27 50.74 74.55 ;
      RECT  49.18 75.27 49.32 74.56 ;
      RECT  50.6 74.41 50.74 69.53 ;
      RECT  50.02 74.63 50.34 74.55 ;
      RECT  49.18 74.56 49.83 74.42 ;
      RECT  50.02 75.59 50.74 75.73 ;
      RECT  49.51 75.51 49.83 75.58 ;
      RECT  49.51 75.72 49.83 75.83 ;
      RECT  50.02 75.73 50.34 75.83 ;
      RECT  49.18 75.72 49.32 80.61 ;
      RECT  50.6 74.87 50.74 75.59 ;
      RECT  49.18 74.87 49.32 75.58 ;
      RECT  50.6 75.73 50.74 80.61 ;
      RECT  50.02 75.51 50.34 75.59 ;
      RECT  49.18 75.58 49.83 75.72 ;
      RECT  50.02 84.73 50.74 84.59 ;
      RECT  49.51 84.81 49.83 84.74 ;
      RECT  49.51 84.6 49.83 84.49 ;
      RECT  50.02 84.59 50.34 84.49 ;
      RECT  49.18 84.6 49.32 79.71 ;
      RECT  50.6 85.45 50.74 84.73 ;
      RECT  49.18 85.45 49.32 84.74 ;
      RECT  50.6 84.59 50.74 79.71 ;
      RECT  50.02 84.81 50.34 84.73 ;
      RECT  49.18 84.74 49.83 84.6 ;
      RECT  50.02 85.77 50.74 85.91 ;
      RECT  49.51 85.69 49.83 85.76 ;
      RECT  49.51 85.9 49.83 86.01 ;
      RECT  50.02 85.91 50.34 86.01 ;
      RECT  49.18 85.9 49.32 90.79 ;
      RECT  50.6 85.05 50.74 85.77 ;
      RECT  49.18 85.05 49.32 85.76 ;
      RECT  50.6 85.91 50.74 90.79 ;
      RECT  50.02 85.69 50.34 85.77 ;
      RECT  49.18 85.76 49.83 85.9 ;
      RECT  50.02 94.91 50.74 94.77 ;
      RECT  49.51 94.99 49.83 94.92 ;
      RECT  49.51 94.78 49.83 94.67 ;
      RECT  50.02 94.77 50.34 94.67 ;
      RECT  49.18 94.78 49.32 89.89 ;
      RECT  50.6 95.63 50.74 94.91 ;
      RECT  49.18 95.63 49.32 94.92 ;
      RECT  50.6 94.77 50.74 89.89 ;
      RECT  50.02 94.99 50.34 94.91 ;
      RECT  49.18 94.92 49.83 94.78 ;
      RECT  50.02 95.95 50.74 96.09 ;
      RECT  49.51 95.87 49.83 95.94 ;
      RECT  49.51 96.08 49.83 96.19 ;
      RECT  50.02 96.09 50.34 96.19 ;
      RECT  49.18 96.08 49.32 100.97 ;
      RECT  50.6 95.23 50.74 95.95 ;
      RECT  49.18 95.23 49.32 95.94 ;
      RECT  50.6 96.09 50.74 100.97 ;
      RECT  50.02 95.87 50.34 95.95 ;
      RECT  49.18 95.94 49.83 96.08 ;
      RECT  50.02 105.09 50.74 104.95 ;
      RECT  49.51 105.17 49.83 105.1 ;
      RECT  49.51 104.96 49.83 104.85 ;
      RECT  50.02 104.95 50.34 104.85 ;
      RECT  49.18 104.96 49.32 100.07 ;
      RECT  50.6 105.81 50.74 105.09 ;
      RECT  49.18 105.81 49.32 105.1 ;
      RECT  50.6 104.95 50.74 100.07 ;
      RECT  50.02 105.17 50.34 105.09 ;
      RECT  49.18 105.1 49.83 104.96 ;
      RECT  50.02 106.13 50.74 106.27 ;
      RECT  49.51 106.05 49.83 106.12 ;
      RECT  49.51 106.26 49.83 106.37 ;
      RECT  50.02 106.27 50.34 106.37 ;
      RECT  49.18 106.26 49.32 111.15 ;
      RECT  50.6 105.41 50.74 106.13 ;
      RECT  49.18 105.41 49.32 106.12 ;
      RECT  50.6 106.27 50.74 111.15 ;
      RECT  50.02 106.05 50.34 106.13 ;
      RECT  49.18 106.12 49.83 106.26 ;
      RECT  50.02 115.27 50.74 115.13 ;
      RECT  49.51 115.35 49.83 115.28 ;
      RECT  49.51 115.14 49.83 115.03 ;
      RECT  50.02 115.13 50.34 115.03 ;
      RECT  49.18 115.14 49.32 110.25 ;
      RECT  50.6 115.99 50.74 115.27 ;
      RECT  49.18 115.99 49.32 115.28 ;
      RECT  50.6 115.13 50.74 110.25 ;
      RECT  50.02 115.35 50.34 115.27 ;
      RECT  49.18 115.28 49.83 115.14 ;
      RECT  52.62 34.87 53.34 35.01 ;
      RECT  52.11 34.79 52.43 34.86 ;
      RECT  52.11 35.0 52.43 35.11 ;
      RECT  52.62 35.01 52.94 35.11 ;
      RECT  51.78 35.0 51.92 39.89 ;
      RECT  53.2 34.15 53.34 34.87 ;
      RECT  51.78 34.15 51.92 34.86 ;
      RECT  53.2 35.01 53.34 39.89 ;
      RECT  52.62 34.79 52.94 34.87 ;
      RECT  51.78 34.86 52.43 35.0 ;
      RECT  52.62 44.01 53.34 43.87 ;
      RECT  52.11 44.09 52.43 44.02 ;
      RECT  52.11 43.88 52.43 43.77 ;
      RECT  52.62 43.87 52.94 43.77 ;
      RECT  51.78 43.88 51.92 38.99 ;
      RECT  53.2 44.73 53.34 44.01 ;
      RECT  51.78 44.73 51.92 44.02 ;
      RECT  53.2 43.87 53.34 38.99 ;
      RECT  52.62 44.09 52.94 44.01 ;
      RECT  51.78 44.02 52.43 43.88 ;
      RECT  52.62 45.05 53.34 45.19 ;
      RECT  52.11 44.97 52.43 45.04 ;
      RECT  52.11 45.18 52.43 45.29 ;
      RECT  52.62 45.19 52.94 45.29 ;
      RECT  51.78 45.18 51.92 50.07 ;
      RECT  53.2 44.33 53.34 45.05 ;
      RECT  51.78 44.33 51.92 45.04 ;
      RECT  53.2 45.19 53.34 50.07 ;
      RECT  52.62 44.97 52.94 45.05 ;
      RECT  51.78 45.04 52.43 45.18 ;
      RECT  52.62 54.19 53.34 54.05 ;
      RECT  52.11 54.27 52.43 54.2 ;
      RECT  52.11 54.06 52.43 53.95 ;
      RECT  52.62 54.05 52.94 53.95 ;
      RECT  51.78 54.06 51.92 49.17 ;
      RECT  53.2 54.91 53.34 54.19 ;
      RECT  51.78 54.91 51.92 54.2 ;
      RECT  53.2 54.05 53.34 49.17 ;
      RECT  52.62 54.27 52.94 54.19 ;
      RECT  51.78 54.2 52.43 54.06 ;
      RECT  52.62 55.23 53.34 55.37 ;
      RECT  52.11 55.15 52.43 55.22 ;
      RECT  52.11 55.36 52.43 55.47 ;
      RECT  52.62 55.37 52.94 55.47 ;
      RECT  51.78 55.36 51.92 60.25 ;
      RECT  53.2 54.51 53.34 55.23 ;
      RECT  51.78 54.51 51.92 55.22 ;
      RECT  53.2 55.37 53.34 60.25 ;
      RECT  52.62 55.15 52.94 55.23 ;
      RECT  51.78 55.22 52.43 55.36 ;
      RECT  52.62 64.37 53.34 64.23 ;
      RECT  52.11 64.45 52.43 64.38 ;
      RECT  52.11 64.24 52.43 64.13 ;
      RECT  52.62 64.23 52.94 64.13 ;
      RECT  51.78 64.24 51.92 59.35 ;
      RECT  53.2 65.09 53.34 64.37 ;
      RECT  51.78 65.09 51.92 64.38 ;
      RECT  53.2 64.23 53.34 59.35 ;
      RECT  52.62 64.45 52.94 64.37 ;
      RECT  51.78 64.38 52.43 64.24 ;
      RECT  52.62 65.41 53.34 65.55 ;
      RECT  52.11 65.33 52.43 65.4 ;
      RECT  52.11 65.54 52.43 65.65 ;
      RECT  52.62 65.55 52.94 65.65 ;
      RECT  51.78 65.54 51.92 70.43 ;
      RECT  53.2 64.69 53.34 65.41 ;
      RECT  51.78 64.69 51.92 65.4 ;
      RECT  53.2 65.55 53.34 70.43 ;
      RECT  52.62 65.33 52.94 65.41 ;
      RECT  51.78 65.4 52.43 65.54 ;
      RECT  52.62 74.55 53.34 74.41 ;
      RECT  52.11 74.63 52.43 74.56 ;
      RECT  52.11 74.42 52.43 74.31 ;
      RECT  52.62 74.41 52.94 74.31 ;
      RECT  51.78 74.42 51.92 69.53 ;
      RECT  53.2 75.27 53.34 74.55 ;
      RECT  51.78 75.27 51.92 74.56 ;
      RECT  53.2 74.41 53.34 69.53 ;
      RECT  52.62 74.63 52.94 74.55 ;
      RECT  51.78 74.56 52.43 74.42 ;
      RECT  52.62 75.59 53.34 75.73 ;
      RECT  52.11 75.51 52.43 75.58 ;
      RECT  52.11 75.72 52.43 75.83 ;
      RECT  52.62 75.73 52.94 75.83 ;
      RECT  51.78 75.72 51.92 80.61 ;
      RECT  53.2 74.87 53.34 75.59 ;
      RECT  51.78 74.87 51.92 75.58 ;
      RECT  53.2 75.73 53.34 80.61 ;
      RECT  52.62 75.51 52.94 75.59 ;
      RECT  51.78 75.58 52.43 75.72 ;
      RECT  52.62 84.73 53.34 84.59 ;
      RECT  52.11 84.81 52.43 84.74 ;
      RECT  52.11 84.6 52.43 84.49 ;
      RECT  52.62 84.59 52.94 84.49 ;
      RECT  51.78 84.6 51.92 79.71 ;
      RECT  53.2 85.45 53.34 84.73 ;
      RECT  51.78 85.45 51.92 84.74 ;
      RECT  53.2 84.59 53.34 79.71 ;
      RECT  52.62 84.81 52.94 84.73 ;
      RECT  51.78 84.74 52.43 84.6 ;
      RECT  52.62 85.77 53.34 85.91 ;
      RECT  52.11 85.69 52.43 85.76 ;
      RECT  52.11 85.9 52.43 86.01 ;
      RECT  52.62 85.91 52.94 86.01 ;
      RECT  51.78 85.9 51.92 90.79 ;
      RECT  53.2 85.05 53.34 85.77 ;
      RECT  51.78 85.05 51.92 85.76 ;
      RECT  53.2 85.91 53.34 90.79 ;
      RECT  52.62 85.69 52.94 85.77 ;
      RECT  51.78 85.76 52.43 85.9 ;
      RECT  52.62 94.91 53.34 94.77 ;
      RECT  52.11 94.99 52.43 94.92 ;
      RECT  52.11 94.78 52.43 94.67 ;
      RECT  52.62 94.77 52.94 94.67 ;
      RECT  51.78 94.78 51.92 89.89 ;
      RECT  53.2 95.63 53.34 94.91 ;
      RECT  51.78 95.63 51.92 94.92 ;
      RECT  53.2 94.77 53.34 89.89 ;
      RECT  52.62 94.99 52.94 94.91 ;
      RECT  51.78 94.92 52.43 94.78 ;
      RECT  52.62 95.95 53.34 96.09 ;
      RECT  52.11 95.87 52.43 95.94 ;
      RECT  52.11 96.08 52.43 96.19 ;
      RECT  52.62 96.09 52.94 96.19 ;
      RECT  51.78 96.08 51.92 100.97 ;
      RECT  53.2 95.23 53.34 95.95 ;
      RECT  51.78 95.23 51.92 95.94 ;
      RECT  53.2 96.09 53.34 100.97 ;
      RECT  52.62 95.87 52.94 95.95 ;
      RECT  51.78 95.94 52.43 96.08 ;
      RECT  52.62 105.09 53.34 104.95 ;
      RECT  52.11 105.17 52.43 105.1 ;
      RECT  52.11 104.96 52.43 104.85 ;
      RECT  52.62 104.95 52.94 104.85 ;
      RECT  51.78 104.96 51.92 100.07 ;
      RECT  53.2 105.81 53.34 105.09 ;
      RECT  51.78 105.81 51.92 105.1 ;
      RECT  53.2 104.95 53.34 100.07 ;
      RECT  52.62 105.17 52.94 105.09 ;
      RECT  51.78 105.1 52.43 104.96 ;
      RECT  52.62 106.13 53.34 106.27 ;
      RECT  52.11 106.05 52.43 106.12 ;
      RECT  52.11 106.26 52.43 106.37 ;
      RECT  52.62 106.27 52.94 106.37 ;
      RECT  51.78 106.26 51.92 111.15 ;
      RECT  53.2 105.41 53.34 106.13 ;
      RECT  51.78 105.41 51.92 106.12 ;
      RECT  53.2 106.27 53.34 111.15 ;
      RECT  52.62 106.05 52.94 106.13 ;
      RECT  51.78 106.12 52.43 106.26 ;
      RECT  52.62 115.27 53.34 115.13 ;
      RECT  52.11 115.35 52.43 115.28 ;
      RECT  52.11 115.14 52.43 115.03 ;
      RECT  52.62 115.13 52.94 115.03 ;
      RECT  51.78 115.14 51.92 110.25 ;
      RECT  53.2 115.99 53.34 115.27 ;
      RECT  51.78 115.99 51.92 115.28 ;
      RECT  53.2 115.13 53.34 110.25 ;
      RECT  52.62 115.35 52.94 115.27 ;
      RECT  51.78 115.28 52.43 115.14 ;
      RECT  49.18 34.35 49.83 115.79 ;
      RECT  50.02 34.35 50.74 115.79 ;
      RECT  51.78 34.35 52.43 115.79 ;
      RECT  52.62 34.35 53.34 115.79 ;
      RECT  47.42 24.69 48.14 24.83 ;
      RECT  46.91 24.61 47.23 24.68 ;
      RECT  46.91 24.82 47.23 24.93 ;
      RECT  47.42 24.83 47.74 24.93 ;
      RECT  46.58 24.82 46.72 29.71 ;
      RECT  48.0 23.97 48.14 24.69 ;
      RECT  46.58 23.97 46.72 24.68 ;
      RECT  48.0 24.83 48.14 29.71 ;
      RECT  47.42 24.61 47.74 24.69 ;
      RECT  46.58 24.68 47.23 24.82 ;
      RECT  47.42 33.83 48.14 33.69 ;
      RECT  46.91 33.91 47.23 33.84 ;
      RECT  46.91 33.7 47.23 33.59 ;
      RECT  47.42 33.69 47.74 33.59 ;
      RECT  46.58 33.7 46.72 28.81 ;
      RECT  48.0 34.55 48.14 33.83 ;
      RECT  46.58 34.55 46.72 33.84 ;
      RECT  48.0 33.69 48.14 28.81 ;
      RECT  47.42 33.91 47.74 33.83 ;
      RECT  46.58 33.84 47.23 33.7 ;
      RECT  47.42 34.87 48.14 35.01 ;
      RECT  46.91 34.79 47.23 34.86 ;
      RECT  46.91 35.0 47.23 35.11 ;
      RECT  47.42 35.01 47.74 35.11 ;
      RECT  46.58 35.0 46.72 39.89 ;
      RECT  48.0 34.15 48.14 34.87 ;
      RECT  46.58 34.15 46.72 34.86 ;
      RECT  48.0 35.01 48.14 39.89 ;
      RECT  47.42 34.79 47.74 34.87 ;
      RECT  46.58 34.86 47.23 35.0 ;
      RECT  47.42 44.01 48.14 43.87 ;
      RECT  46.91 44.09 47.23 44.02 ;
      RECT  46.91 43.88 47.23 43.77 ;
      RECT  47.42 43.87 47.74 43.77 ;
      RECT  46.58 43.88 46.72 38.99 ;
      RECT  48.0 44.73 48.14 44.01 ;
      RECT  46.58 44.73 46.72 44.02 ;
      RECT  48.0 43.87 48.14 38.99 ;
      RECT  47.42 44.09 47.74 44.01 ;
      RECT  46.58 44.02 47.23 43.88 ;
      RECT  47.42 45.05 48.14 45.19 ;
      RECT  46.91 44.97 47.23 45.04 ;
      RECT  46.91 45.18 47.23 45.29 ;
      RECT  47.42 45.19 47.74 45.29 ;
      RECT  46.58 45.18 46.72 50.07 ;
      RECT  48.0 44.33 48.14 45.05 ;
      RECT  46.58 44.33 46.72 45.04 ;
      RECT  48.0 45.19 48.14 50.07 ;
      RECT  47.42 44.97 47.74 45.05 ;
      RECT  46.58 45.04 47.23 45.18 ;
      RECT  47.42 54.19 48.14 54.05 ;
      RECT  46.91 54.27 47.23 54.2 ;
      RECT  46.91 54.06 47.23 53.95 ;
      RECT  47.42 54.05 47.74 53.95 ;
      RECT  46.58 54.06 46.72 49.17 ;
      RECT  48.0 54.91 48.14 54.19 ;
      RECT  46.58 54.91 46.72 54.2 ;
      RECT  48.0 54.05 48.14 49.17 ;
      RECT  47.42 54.27 47.74 54.19 ;
      RECT  46.58 54.2 47.23 54.06 ;
      RECT  47.42 55.23 48.14 55.37 ;
      RECT  46.91 55.15 47.23 55.22 ;
      RECT  46.91 55.36 47.23 55.47 ;
      RECT  47.42 55.37 47.74 55.47 ;
      RECT  46.58 55.36 46.72 60.25 ;
      RECT  48.0 54.51 48.14 55.23 ;
      RECT  46.58 54.51 46.72 55.22 ;
      RECT  48.0 55.37 48.14 60.25 ;
      RECT  47.42 55.15 47.74 55.23 ;
      RECT  46.58 55.22 47.23 55.36 ;
      RECT  47.42 64.37 48.14 64.23 ;
      RECT  46.91 64.45 47.23 64.38 ;
      RECT  46.91 64.24 47.23 64.13 ;
      RECT  47.42 64.23 47.74 64.13 ;
      RECT  46.58 64.24 46.72 59.35 ;
      RECT  48.0 65.09 48.14 64.37 ;
      RECT  46.58 65.09 46.72 64.38 ;
      RECT  48.0 64.23 48.14 59.35 ;
      RECT  47.42 64.45 47.74 64.37 ;
      RECT  46.58 64.38 47.23 64.24 ;
      RECT  47.42 65.41 48.14 65.55 ;
      RECT  46.91 65.33 47.23 65.4 ;
      RECT  46.91 65.54 47.23 65.65 ;
      RECT  47.42 65.55 47.74 65.65 ;
      RECT  46.58 65.54 46.72 70.43 ;
      RECT  48.0 64.69 48.14 65.41 ;
      RECT  46.58 64.69 46.72 65.4 ;
      RECT  48.0 65.55 48.14 70.43 ;
      RECT  47.42 65.33 47.74 65.41 ;
      RECT  46.58 65.4 47.23 65.54 ;
      RECT  47.42 74.55 48.14 74.41 ;
      RECT  46.91 74.63 47.23 74.56 ;
      RECT  46.91 74.42 47.23 74.31 ;
      RECT  47.42 74.41 47.74 74.31 ;
      RECT  46.58 74.42 46.72 69.53 ;
      RECT  48.0 75.27 48.14 74.55 ;
      RECT  46.58 75.27 46.72 74.56 ;
      RECT  48.0 74.41 48.14 69.53 ;
      RECT  47.42 74.63 47.74 74.55 ;
      RECT  46.58 74.56 47.23 74.42 ;
      RECT  47.42 75.59 48.14 75.73 ;
      RECT  46.91 75.51 47.23 75.58 ;
      RECT  46.91 75.72 47.23 75.83 ;
      RECT  47.42 75.73 47.74 75.83 ;
      RECT  46.58 75.72 46.72 80.61 ;
      RECT  48.0 74.87 48.14 75.59 ;
      RECT  46.58 74.87 46.72 75.58 ;
      RECT  48.0 75.73 48.14 80.61 ;
      RECT  47.42 75.51 47.74 75.59 ;
      RECT  46.58 75.58 47.23 75.72 ;
      RECT  47.42 84.73 48.14 84.59 ;
      RECT  46.91 84.81 47.23 84.74 ;
      RECT  46.91 84.6 47.23 84.49 ;
      RECT  47.42 84.59 47.74 84.49 ;
      RECT  46.58 84.6 46.72 79.71 ;
      RECT  48.0 85.45 48.14 84.73 ;
      RECT  46.58 85.45 46.72 84.74 ;
      RECT  48.0 84.59 48.14 79.71 ;
      RECT  47.42 84.81 47.74 84.73 ;
      RECT  46.58 84.74 47.23 84.6 ;
      RECT  47.42 85.77 48.14 85.91 ;
      RECT  46.91 85.69 47.23 85.76 ;
      RECT  46.91 85.9 47.23 86.01 ;
      RECT  47.42 85.91 47.74 86.01 ;
      RECT  46.58 85.9 46.72 90.79 ;
      RECT  48.0 85.05 48.14 85.77 ;
      RECT  46.58 85.05 46.72 85.76 ;
      RECT  48.0 85.91 48.14 90.79 ;
      RECT  47.42 85.69 47.74 85.77 ;
      RECT  46.58 85.76 47.23 85.9 ;
      RECT  47.42 94.91 48.14 94.77 ;
      RECT  46.91 94.99 47.23 94.92 ;
      RECT  46.91 94.78 47.23 94.67 ;
      RECT  47.42 94.77 47.74 94.67 ;
      RECT  46.58 94.78 46.72 89.89 ;
      RECT  48.0 95.63 48.14 94.91 ;
      RECT  46.58 95.63 46.72 94.92 ;
      RECT  48.0 94.77 48.14 89.89 ;
      RECT  47.42 94.99 47.74 94.91 ;
      RECT  46.58 94.92 47.23 94.78 ;
      RECT  47.42 95.95 48.14 96.09 ;
      RECT  46.91 95.87 47.23 95.94 ;
      RECT  46.91 96.08 47.23 96.19 ;
      RECT  47.42 96.09 47.74 96.19 ;
      RECT  46.58 96.08 46.72 100.97 ;
      RECT  48.0 95.23 48.14 95.95 ;
      RECT  46.58 95.23 46.72 95.94 ;
      RECT  48.0 96.09 48.14 100.97 ;
      RECT  47.42 95.87 47.74 95.95 ;
      RECT  46.58 95.94 47.23 96.08 ;
      RECT  47.42 105.09 48.14 104.95 ;
      RECT  46.91 105.17 47.23 105.1 ;
      RECT  46.91 104.96 47.23 104.85 ;
      RECT  47.42 104.95 47.74 104.85 ;
      RECT  46.58 104.96 46.72 100.07 ;
      RECT  48.0 105.81 48.14 105.09 ;
      RECT  46.58 105.81 46.72 105.1 ;
      RECT  48.0 104.95 48.14 100.07 ;
      RECT  47.42 105.17 47.74 105.09 ;
      RECT  46.58 105.1 47.23 104.96 ;
      RECT  47.42 106.13 48.14 106.27 ;
      RECT  46.91 106.05 47.23 106.12 ;
      RECT  46.91 106.26 47.23 106.37 ;
      RECT  47.42 106.27 47.74 106.37 ;
      RECT  46.58 106.26 46.72 111.15 ;
      RECT  48.0 105.41 48.14 106.13 ;
      RECT  46.58 105.41 46.72 106.12 ;
      RECT  48.0 106.27 48.14 111.15 ;
      RECT  47.42 106.05 47.74 106.13 ;
      RECT  46.58 106.12 47.23 106.26 ;
      RECT  47.42 115.27 48.14 115.13 ;
      RECT  46.91 115.35 47.23 115.28 ;
      RECT  46.91 115.14 47.23 115.03 ;
      RECT  47.42 115.13 47.74 115.03 ;
      RECT  46.58 115.14 46.72 110.25 ;
      RECT  48.0 115.99 48.14 115.27 ;
      RECT  46.58 115.99 46.72 115.28 ;
      RECT  48.0 115.13 48.14 110.25 ;
      RECT  47.42 115.35 47.74 115.27 ;
      RECT  46.58 115.28 47.23 115.14 ;
      RECT  47.42 116.31 48.14 116.45 ;
      RECT  46.91 116.23 47.23 116.3 ;
      RECT  46.91 116.44 47.23 116.55 ;
      RECT  47.42 116.45 47.74 116.55 ;
      RECT  46.58 116.44 46.72 121.33 ;
      RECT  48.0 115.59 48.14 116.31 ;
      RECT  46.58 115.59 46.72 116.3 ;
      RECT  48.0 116.45 48.14 121.33 ;
      RECT  47.42 116.23 47.74 116.31 ;
      RECT  46.58 116.3 47.23 116.44 ;
      RECT  46.58 24.17 47.23 120.88 ;
      RECT  47.42 24.17 48.14 120.88 ;
      RECT  50.02 33.83 50.74 33.69 ;
      RECT  49.51 33.91 49.83 33.84 ;
      RECT  49.51 33.7 49.83 33.59 ;
      RECT  50.02 33.69 50.34 33.59 ;
      RECT  49.18 33.7 49.32 28.81 ;
      RECT  50.6 34.55 50.74 33.83 ;
      RECT  49.18 34.55 49.32 33.84 ;
      RECT  50.6 33.69 50.74 28.81 ;
      RECT  50.02 33.91 50.34 33.83 ;
      RECT  49.18 33.84 49.83 33.7 ;
      RECT  52.62 33.83 53.34 33.69 ;
      RECT  52.11 33.91 52.43 33.84 ;
      RECT  52.11 33.7 52.43 33.59 ;
      RECT  52.62 33.69 52.94 33.59 ;
      RECT  51.78 33.7 51.92 28.81 ;
      RECT  53.2 34.55 53.34 33.83 ;
      RECT  51.78 34.55 51.92 33.84 ;
      RECT  53.2 33.69 53.34 28.81 ;
      RECT  52.62 33.91 52.94 33.83 ;
      RECT  51.78 33.84 52.43 33.7 ;
      RECT  49.18 34.35 49.83 29.26 ;
      RECT  50.02 34.35 50.74 29.26 ;
      RECT  51.78 34.35 52.43 29.26 ;
      RECT  52.62 34.35 53.34 29.26 ;
      RECT  50.02 24.69 50.74 24.83 ;
      RECT  49.51 24.61 49.83 24.68 ;
      RECT  49.51 24.82 49.83 24.93 ;
      RECT  50.02 24.83 50.34 24.93 ;
      RECT  49.18 24.82 49.32 29.71 ;
      RECT  50.6 23.97 50.74 24.69 ;
      RECT  49.18 23.97 49.32 24.68 ;
      RECT  50.6 24.83 50.74 29.71 ;
      RECT  50.02 24.61 50.34 24.69 ;
      RECT  49.18 24.68 49.83 24.82 ;
      RECT  52.62 24.69 53.34 24.83 ;
      RECT  52.11 24.61 52.43 24.68 ;
      RECT  52.11 24.82 52.43 24.93 ;
      RECT  52.62 24.83 52.94 24.93 ;
      RECT  51.78 24.82 51.92 29.71 ;
      RECT  53.2 23.97 53.34 24.69 ;
      RECT  51.78 23.97 51.92 24.68 ;
      RECT  53.2 24.83 53.34 29.71 ;
      RECT  52.62 24.61 52.94 24.69 ;
      RECT  51.78 24.68 52.43 24.82 ;
      RECT  49.18 24.17 49.83 29.26 ;
      RECT  50.02 24.17 50.74 29.26 ;
      RECT  51.78 24.17 52.43 29.26 ;
      RECT  52.62 24.17 53.34 29.26 ;
      RECT  50.02 116.31 50.74 116.45 ;
      RECT  49.51 116.23 49.83 116.3 ;
      RECT  49.51 116.44 49.83 116.55 ;
      RECT  50.02 116.45 50.34 116.55 ;
      RECT  49.18 116.44 49.32 121.33 ;
      RECT  50.6 115.59 50.74 116.31 ;
      RECT  49.18 115.59 49.32 116.3 ;
      RECT  50.6 116.45 50.74 121.33 ;
      RECT  50.02 116.23 50.34 116.31 ;
      RECT  49.18 116.3 49.83 116.44 ;
      RECT  52.62 116.31 53.34 116.45 ;
      RECT  52.11 116.23 52.43 116.3 ;
      RECT  52.11 116.44 52.43 116.55 ;
      RECT  52.62 116.45 52.94 116.55 ;
      RECT  51.78 116.44 51.92 121.33 ;
      RECT  53.2 115.59 53.34 116.31 ;
      RECT  51.78 115.59 51.92 116.3 ;
      RECT  53.2 116.45 53.34 121.33 ;
      RECT  52.62 116.23 52.94 116.31 ;
      RECT  51.78 116.3 52.43 116.44 ;
      RECT  49.18 115.79 49.83 120.88 ;
      RECT  50.02 115.79 50.74 120.88 ;
      RECT  51.78 115.79 52.43 120.88 ;
      RECT  52.62 115.79 53.34 120.88 ;
      RECT  44.82 24.69 45.54 24.83 ;
      RECT  44.31 24.61 44.63 24.68 ;
      RECT  44.31 24.82 44.63 24.93 ;
      RECT  44.82 24.83 45.14 24.93 ;
      RECT  43.98 24.82 44.12 29.71 ;
      RECT  45.4 23.97 45.54 24.69 ;
      RECT  43.98 23.97 44.12 24.68 ;
      RECT  45.4 24.83 45.54 29.71 ;
      RECT  44.82 24.61 45.14 24.69 ;
      RECT  43.98 24.68 44.63 24.82 ;
      RECT  44.82 33.83 45.54 33.69 ;
      RECT  44.31 33.91 44.63 33.84 ;
      RECT  44.31 33.7 44.63 33.59 ;
      RECT  44.82 33.69 45.14 33.59 ;
      RECT  43.98 33.7 44.12 28.81 ;
      RECT  45.4 34.55 45.54 33.83 ;
      RECT  43.98 34.55 44.12 33.84 ;
      RECT  45.4 33.69 45.54 28.81 ;
      RECT  44.82 33.91 45.14 33.83 ;
      RECT  43.98 33.84 44.63 33.7 ;
      RECT  44.82 34.87 45.54 35.01 ;
      RECT  44.31 34.79 44.63 34.86 ;
      RECT  44.31 35.0 44.63 35.11 ;
      RECT  44.82 35.01 45.14 35.11 ;
      RECT  43.98 35.0 44.12 39.89 ;
      RECT  45.4 34.15 45.54 34.87 ;
      RECT  43.98 34.15 44.12 34.86 ;
      RECT  45.4 35.01 45.54 39.89 ;
      RECT  44.82 34.79 45.14 34.87 ;
      RECT  43.98 34.86 44.63 35.0 ;
      RECT  44.82 44.01 45.54 43.87 ;
      RECT  44.31 44.09 44.63 44.02 ;
      RECT  44.31 43.88 44.63 43.77 ;
      RECT  44.82 43.87 45.14 43.77 ;
      RECT  43.98 43.88 44.12 38.99 ;
      RECT  45.4 44.73 45.54 44.01 ;
      RECT  43.98 44.73 44.12 44.02 ;
      RECT  45.4 43.87 45.54 38.99 ;
      RECT  44.82 44.09 45.14 44.01 ;
      RECT  43.98 44.02 44.63 43.88 ;
      RECT  44.82 45.05 45.54 45.19 ;
      RECT  44.31 44.97 44.63 45.04 ;
      RECT  44.31 45.18 44.63 45.29 ;
      RECT  44.82 45.19 45.14 45.29 ;
      RECT  43.98 45.18 44.12 50.07 ;
      RECT  45.4 44.33 45.54 45.05 ;
      RECT  43.98 44.33 44.12 45.04 ;
      RECT  45.4 45.19 45.54 50.07 ;
      RECT  44.82 44.97 45.14 45.05 ;
      RECT  43.98 45.04 44.63 45.18 ;
      RECT  44.82 54.19 45.54 54.05 ;
      RECT  44.31 54.27 44.63 54.2 ;
      RECT  44.31 54.06 44.63 53.95 ;
      RECT  44.82 54.05 45.14 53.95 ;
      RECT  43.98 54.06 44.12 49.17 ;
      RECT  45.4 54.91 45.54 54.19 ;
      RECT  43.98 54.91 44.12 54.2 ;
      RECT  45.4 54.05 45.54 49.17 ;
      RECT  44.82 54.27 45.14 54.19 ;
      RECT  43.98 54.2 44.63 54.06 ;
      RECT  44.82 55.23 45.54 55.37 ;
      RECT  44.31 55.15 44.63 55.22 ;
      RECT  44.31 55.36 44.63 55.47 ;
      RECT  44.82 55.37 45.14 55.47 ;
      RECT  43.98 55.36 44.12 60.25 ;
      RECT  45.4 54.51 45.54 55.23 ;
      RECT  43.98 54.51 44.12 55.22 ;
      RECT  45.4 55.37 45.54 60.25 ;
      RECT  44.82 55.15 45.14 55.23 ;
      RECT  43.98 55.22 44.63 55.36 ;
      RECT  44.82 64.37 45.54 64.23 ;
      RECT  44.31 64.45 44.63 64.38 ;
      RECT  44.31 64.24 44.63 64.13 ;
      RECT  44.82 64.23 45.14 64.13 ;
      RECT  43.98 64.24 44.12 59.35 ;
      RECT  45.4 65.09 45.54 64.37 ;
      RECT  43.98 65.09 44.12 64.38 ;
      RECT  45.4 64.23 45.54 59.35 ;
      RECT  44.82 64.45 45.14 64.37 ;
      RECT  43.98 64.38 44.63 64.24 ;
      RECT  44.82 65.41 45.54 65.55 ;
      RECT  44.31 65.33 44.63 65.4 ;
      RECT  44.31 65.54 44.63 65.65 ;
      RECT  44.82 65.55 45.14 65.65 ;
      RECT  43.98 65.54 44.12 70.43 ;
      RECT  45.4 64.69 45.54 65.41 ;
      RECT  43.98 64.69 44.12 65.4 ;
      RECT  45.4 65.55 45.54 70.43 ;
      RECT  44.82 65.33 45.14 65.41 ;
      RECT  43.98 65.4 44.63 65.54 ;
      RECT  44.82 74.55 45.54 74.41 ;
      RECT  44.31 74.63 44.63 74.56 ;
      RECT  44.31 74.42 44.63 74.31 ;
      RECT  44.82 74.41 45.14 74.31 ;
      RECT  43.98 74.42 44.12 69.53 ;
      RECT  45.4 75.27 45.54 74.55 ;
      RECT  43.98 75.27 44.12 74.56 ;
      RECT  45.4 74.41 45.54 69.53 ;
      RECT  44.82 74.63 45.14 74.55 ;
      RECT  43.98 74.56 44.63 74.42 ;
      RECT  44.82 75.59 45.54 75.73 ;
      RECT  44.31 75.51 44.63 75.58 ;
      RECT  44.31 75.72 44.63 75.83 ;
      RECT  44.82 75.73 45.14 75.83 ;
      RECT  43.98 75.72 44.12 80.61 ;
      RECT  45.4 74.87 45.54 75.59 ;
      RECT  43.98 74.87 44.12 75.58 ;
      RECT  45.4 75.73 45.54 80.61 ;
      RECT  44.82 75.51 45.14 75.59 ;
      RECT  43.98 75.58 44.63 75.72 ;
      RECT  44.82 84.73 45.54 84.59 ;
      RECT  44.31 84.81 44.63 84.74 ;
      RECT  44.31 84.6 44.63 84.49 ;
      RECT  44.82 84.59 45.14 84.49 ;
      RECT  43.98 84.6 44.12 79.71 ;
      RECT  45.4 85.45 45.54 84.73 ;
      RECT  43.98 85.45 44.12 84.74 ;
      RECT  45.4 84.59 45.54 79.71 ;
      RECT  44.82 84.81 45.14 84.73 ;
      RECT  43.98 84.74 44.63 84.6 ;
      RECT  44.82 85.77 45.54 85.91 ;
      RECT  44.31 85.69 44.63 85.76 ;
      RECT  44.31 85.9 44.63 86.01 ;
      RECT  44.82 85.91 45.14 86.01 ;
      RECT  43.98 85.9 44.12 90.79 ;
      RECT  45.4 85.05 45.54 85.77 ;
      RECT  43.98 85.05 44.12 85.76 ;
      RECT  45.4 85.91 45.54 90.79 ;
      RECT  44.82 85.69 45.14 85.77 ;
      RECT  43.98 85.76 44.63 85.9 ;
      RECT  44.82 94.91 45.54 94.77 ;
      RECT  44.31 94.99 44.63 94.92 ;
      RECT  44.31 94.78 44.63 94.67 ;
      RECT  44.82 94.77 45.14 94.67 ;
      RECT  43.98 94.78 44.12 89.89 ;
      RECT  45.4 95.63 45.54 94.91 ;
      RECT  43.98 95.63 44.12 94.92 ;
      RECT  45.4 94.77 45.54 89.89 ;
      RECT  44.82 94.99 45.14 94.91 ;
      RECT  43.98 94.92 44.63 94.78 ;
      RECT  44.82 95.95 45.54 96.09 ;
      RECT  44.31 95.87 44.63 95.94 ;
      RECT  44.31 96.08 44.63 96.19 ;
      RECT  44.82 96.09 45.14 96.19 ;
      RECT  43.98 96.08 44.12 100.97 ;
      RECT  45.4 95.23 45.54 95.95 ;
      RECT  43.98 95.23 44.12 95.94 ;
      RECT  45.4 96.09 45.54 100.97 ;
      RECT  44.82 95.87 45.14 95.95 ;
      RECT  43.98 95.94 44.63 96.08 ;
      RECT  44.82 105.09 45.54 104.95 ;
      RECT  44.31 105.17 44.63 105.1 ;
      RECT  44.31 104.96 44.63 104.85 ;
      RECT  44.82 104.95 45.14 104.85 ;
      RECT  43.98 104.96 44.12 100.07 ;
      RECT  45.4 105.81 45.54 105.09 ;
      RECT  43.98 105.81 44.12 105.1 ;
      RECT  45.4 104.95 45.54 100.07 ;
      RECT  44.82 105.17 45.14 105.09 ;
      RECT  43.98 105.1 44.63 104.96 ;
      RECT  44.82 106.13 45.54 106.27 ;
      RECT  44.31 106.05 44.63 106.12 ;
      RECT  44.31 106.26 44.63 106.37 ;
      RECT  44.82 106.27 45.14 106.37 ;
      RECT  43.98 106.26 44.12 111.15 ;
      RECT  45.4 105.41 45.54 106.13 ;
      RECT  43.98 105.41 44.12 106.12 ;
      RECT  45.4 106.27 45.54 111.15 ;
      RECT  44.82 106.05 45.14 106.13 ;
      RECT  43.98 106.12 44.63 106.26 ;
      RECT  44.82 115.27 45.54 115.13 ;
      RECT  44.31 115.35 44.63 115.28 ;
      RECT  44.31 115.14 44.63 115.03 ;
      RECT  44.82 115.13 45.14 115.03 ;
      RECT  43.98 115.14 44.12 110.25 ;
      RECT  45.4 115.99 45.54 115.27 ;
      RECT  43.98 115.99 44.12 115.28 ;
      RECT  45.4 115.13 45.54 110.25 ;
      RECT  44.82 115.35 45.14 115.27 ;
      RECT  43.98 115.28 44.63 115.14 ;
      RECT  44.82 116.31 45.54 116.45 ;
      RECT  44.31 116.23 44.63 116.3 ;
      RECT  44.31 116.44 44.63 116.55 ;
      RECT  44.82 116.45 45.14 116.55 ;
      RECT  43.98 116.44 44.12 121.33 ;
      RECT  45.4 115.59 45.54 116.31 ;
      RECT  43.98 115.59 44.12 116.3 ;
      RECT  45.4 116.45 45.54 121.33 ;
      RECT  44.82 116.23 45.14 116.31 ;
      RECT  43.98 116.3 44.63 116.44 ;
      RECT  43.98 24.17 44.63 120.88 ;
      RECT  44.82 24.17 45.54 120.88 ;
      RECT  55.22 24.69 55.94 24.83 ;
      RECT  54.71 24.61 55.03 24.68 ;
      RECT  54.71 24.82 55.03 24.93 ;
      RECT  55.22 24.83 55.54 24.93 ;
      RECT  54.38 24.82 54.52 29.71 ;
      RECT  55.8 23.97 55.94 24.69 ;
      RECT  54.38 23.97 54.52 24.68 ;
      RECT  55.8 24.83 55.94 29.71 ;
      RECT  55.22 24.61 55.54 24.69 ;
      RECT  54.38 24.68 55.03 24.82 ;
      RECT  55.22 33.83 55.94 33.69 ;
      RECT  54.71 33.91 55.03 33.84 ;
      RECT  54.71 33.7 55.03 33.59 ;
      RECT  55.22 33.69 55.54 33.59 ;
      RECT  54.38 33.7 54.52 28.81 ;
      RECT  55.8 34.55 55.94 33.83 ;
      RECT  54.38 34.55 54.52 33.84 ;
      RECT  55.8 33.69 55.94 28.81 ;
      RECT  55.22 33.91 55.54 33.83 ;
      RECT  54.38 33.84 55.03 33.7 ;
      RECT  55.22 34.87 55.94 35.01 ;
      RECT  54.71 34.79 55.03 34.86 ;
      RECT  54.71 35.0 55.03 35.11 ;
      RECT  55.22 35.01 55.54 35.11 ;
      RECT  54.38 35.0 54.52 39.89 ;
      RECT  55.8 34.15 55.94 34.87 ;
      RECT  54.38 34.15 54.52 34.86 ;
      RECT  55.8 35.01 55.94 39.89 ;
      RECT  55.22 34.79 55.54 34.87 ;
      RECT  54.38 34.86 55.03 35.0 ;
      RECT  55.22 44.01 55.94 43.87 ;
      RECT  54.71 44.09 55.03 44.02 ;
      RECT  54.71 43.88 55.03 43.77 ;
      RECT  55.22 43.87 55.54 43.77 ;
      RECT  54.38 43.88 54.52 38.99 ;
      RECT  55.8 44.73 55.94 44.01 ;
      RECT  54.38 44.73 54.52 44.02 ;
      RECT  55.8 43.87 55.94 38.99 ;
      RECT  55.22 44.09 55.54 44.01 ;
      RECT  54.38 44.02 55.03 43.88 ;
      RECT  55.22 45.05 55.94 45.19 ;
      RECT  54.71 44.97 55.03 45.04 ;
      RECT  54.71 45.18 55.03 45.29 ;
      RECT  55.22 45.19 55.54 45.29 ;
      RECT  54.38 45.18 54.52 50.07 ;
      RECT  55.8 44.33 55.94 45.05 ;
      RECT  54.38 44.33 54.52 45.04 ;
      RECT  55.8 45.19 55.94 50.07 ;
      RECT  55.22 44.97 55.54 45.05 ;
      RECT  54.38 45.04 55.03 45.18 ;
      RECT  55.22 54.19 55.94 54.05 ;
      RECT  54.71 54.27 55.03 54.2 ;
      RECT  54.71 54.06 55.03 53.95 ;
      RECT  55.22 54.05 55.54 53.95 ;
      RECT  54.38 54.06 54.52 49.17 ;
      RECT  55.8 54.91 55.94 54.19 ;
      RECT  54.38 54.91 54.52 54.2 ;
      RECT  55.8 54.05 55.94 49.17 ;
      RECT  55.22 54.27 55.54 54.19 ;
      RECT  54.38 54.2 55.03 54.06 ;
      RECT  55.22 55.23 55.94 55.37 ;
      RECT  54.71 55.15 55.03 55.22 ;
      RECT  54.71 55.36 55.03 55.47 ;
      RECT  55.22 55.37 55.54 55.47 ;
      RECT  54.38 55.36 54.52 60.25 ;
      RECT  55.8 54.51 55.94 55.23 ;
      RECT  54.38 54.51 54.52 55.22 ;
      RECT  55.8 55.37 55.94 60.25 ;
      RECT  55.22 55.15 55.54 55.23 ;
      RECT  54.38 55.22 55.03 55.36 ;
      RECT  55.22 64.37 55.94 64.23 ;
      RECT  54.71 64.45 55.03 64.38 ;
      RECT  54.71 64.24 55.03 64.13 ;
      RECT  55.22 64.23 55.54 64.13 ;
      RECT  54.38 64.24 54.52 59.35 ;
      RECT  55.8 65.09 55.94 64.37 ;
      RECT  54.38 65.09 54.52 64.38 ;
      RECT  55.8 64.23 55.94 59.35 ;
      RECT  55.22 64.45 55.54 64.37 ;
      RECT  54.38 64.38 55.03 64.24 ;
      RECT  55.22 65.41 55.94 65.55 ;
      RECT  54.71 65.33 55.03 65.4 ;
      RECT  54.71 65.54 55.03 65.65 ;
      RECT  55.22 65.55 55.54 65.65 ;
      RECT  54.38 65.54 54.52 70.43 ;
      RECT  55.8 64.69 55.94 65.41 ;
      RECT  54.38 64.69 54.52 65.4 ;
      RECT  55.8 65.55 55.94 70.43 ;
      RECT  55.22 65.33 55.54 65.41 ;
      RECT  54.38 65.4 55.03 65.54 ;
      RECT  55.22 74.55 55.94 74.41 ;
      RECT  54.71 74.63 55.03 74.56 ;
      RECT  54.71 74.42 55.03 74.31 ;
      RECT  55.22 74.41 55.54 74.31 ;
      RECT  54.38 74.42 54.52 69.53 ;
      RECT  55.8 75.27 55.94 74.55 ;
      RECT  54.38 75.27 54.52 74.56 ;
      RECT  55.8 74.41 55.94 69.53 ;
      RECT  55.22 74.63 55.54 74.55 ;
      RECT  54.38 74.56 55.03 74.42 ;
      RECT  55.22 75.59 55.94 75.73 ;
      RECT  54.71 75.51 55.03 75.58 ;
      RECT  54.71 75.72 55.03 75.83 ;
      RECT  55.22 75.73 55.54 75.83 ;
      RECT  54.38 75.72 54.52 80.61 ;
      RECT  55.8 74.87 55.94 75.59 ;
      RECT  54.38 74.87 54.52 75.58 ;
      RECT  55.8 75.73 55.94 80.61 ;
      RECT  55.22 75.51 55.54 75.59 ;
      RECT  54.38 75.58 55.03 75.72 ;
      RECT  55.22 84.73 55.94 84.59 ;
      RECT  54.71 84.81 55.03 84.74 ;
      RECT  54.71 84.6 55.03 84.49 ;
      RECT  55.22 84.59 55.54 84.49 ;
      RECT  54.38 84.6 54.52 79.71 ;
      RECT  55.8 85.45 55.94 84.73 ;
      RECT  54.38 85.45 54.52 84.74 ;
      RECT  55.8 84.59 55.94 79.71 ;
      RECT  55.22 84.81 55.54 84.73 ;
      RECT  54.38 84.74 55.03 84.6 ;
      RECT  55.22 85.77 55.94 85.91 ;
      RECT  54.71 85.69 55.03 85.76 ;
      RECT  54.71 85.9 55.03 86.01 ;
      RECT  55.22 85.91 55.54 86.01 ;
      RECT  54.38 85.9 54.52 90.79 ;
      RECT  55.8 85.05 55.94 85.77 ;
      RECT  54.38 85.05 54.52 85.76 ;
      RECT  55.8 85.91 55.94 90.79 ;
      RECT  55.22 85.69 55.54 85.77 ;
      RECT  54.38 85.76 55.03 85.9 ;
      RECT  55.22 94.91 55.94 94.77 ;
      RECT  54.71 94.99 55.03 94.92 ;
      RECT  54.71 94.78 55.03 94.67 ;
      RECT  55.22 94.77 55.54 94.67 ;
      RECT  54.38 94.78 54.52 89.89 ;
      RECT  55.8 95.63 55.94 94.91 ;
      RECT  54.38 95.63 54.52 94.92 ;
      RECT  55.8 94.77 55.94 89.89 ;
      RECT  55.22 94.99 55.54 94.91 ;
      RECT  54.38 94.92 55.03 94.78 ;
      RECT  55.22 95.95 55.94 96.09 ;
      RECT  54.71 95.87 55.03 95.94 ;
      RECT  54.71 96.08 55.03 96.19 ;
      RECT  55.22 96.09 55.54 96.19 ;
      RECT  54.38 96.08 54.52 100.97 ;
      RECT  55.8 95.23 55.94 95.95 ;
      RECT  54.38 95.23 54.52 95.94 ;
      RECT  55.8 96.09 55.94 100.97 ;
      RECT  55.22 95.87 55.54 95.95 ;
      RECT  54.38 95.94 55.03 96.08 ;
      RECT  55.22 105.09 55.94 104.95 ;
      RECT  54.71 105.17 55.03 105.1 ;
      RECT  54.71 104.96 55.03 104.85 ;
      RECT  55.22 104.95 55.54 104.85 ;
      RECT  54.38 104.96 54.52 100.07 ;
      RECT  55.8 105.81 55.94 105.09 ;
      RECT  54.38 105.81 54.52 105.1 ;
      RECT  55.8 104.95 55.94 100.07 ;
      RECT  55.22 105.17 55.54 105.09 ;
      RECT  54.38 105.1 55.03 104.96 ;
      RECT  55.22 106.13 55.94 106.27 ;
      RECT  54.71 106.05 55.03 106.12 ;
      RECT  54.71 106.26 55.03 106.37 ;
      RECT  55.22 106.27 55.54 106.37 ;
      RECT  54.38 106.26 54.52 111.15 ;
      RECT  55.8 105.41 55.94 106.13 ;
      RECT  54.38 105.41 54.52 106.12 ;
      RECT  55.8 106.27 55.94 111.15 ;
      RECT  55.22 106.05 55.54 106.13 ;
      RECT  54.38 106.12 55.03 106.26 ;
      RECT  55.22 115.27 55.94 115.13 ;
      RECT  54.71 115.35 55.03 115.28 ;
      RECT  54.71 115.14 55.03 115.03 ;
      RECT  55.22 115.13 55.54 115.03 ;
      RECT  54.38 115.14 54.52 110.25 ;
      RECT  55.8 115.99 55.94 115.27 ;
      RECT  54.38 115.99 54.52 115.28 ;
      RECT  55.8 115.13 55.94 110.25 ;
      RECT  55.22 115.35 55.54 115.27 ;
      RECT  54.38 115.28 55.03 115.14 ;
      RECT  55.22 116.31 55.94 116.45 ;
      RECT  54.71 116.23 55.03 116.3 ;
      RECT  54.71 116.44 55.03 116.55 ;
      RECT  55.22 116.45 55.54 116.55 ;
      RECT  54.38 116.44 54.52 121.33 ;
      RECT  55.8 115.59 55.94 116.31 ;
      RECT  54.38 115.59 54.52 116.3 ;
      RECT  55.8 116.45 55.94 121.33 ;
      RECT  55.22 116.23 55.54 116.31 ;
      RECT  54.38 116.3 55.03 116.44 ;
      RECT  54.38 24.17 55.03 120.88 ;
      RECT  55.22 24.17 55.94 120.88 ;
      RECT  46.58 24.17 47.23 120.88 ;
      RECT  47.42 24.17 48.14 120.88 ;
      RECT  49.18 24.17 49.83 120.88 ;
      RECT  50.02 24.17 50.74 120.88 ;
      RECT  51.78 24.17 52.43 120.88 ;
      RECT  52.62 24.17 53.34 120.88 ;
      RECT  46.64 15.19 46.78 22.19 ;
      RECT  47.92 15.19 48.06 22.19 ;
      RECT  49.24 15.19 49.38 22.19 ;
      RECT  50.52 15.19 50.66 22.19 ;
      RECT  51.84 15.19 51.98 22.19 ;
      RECT  53.12 15.19 53.26 22.19 ;
      RECT  46.64 15.19 46.78 22.19 ;
      RECT  47.92 15.19 48.06 22.19 ;
      RECT  49.24 15.19 49.38 22.19 ;
      RECT  50.52 15.19 50.66 22.19 ;
      RECT  51.84 15.19 51.98 22.19 ;
      RECT  53.12 15.19 53.26 22.19 ;
      RECT  48.36 8.63 48.69 13.67 ;
      RECT  53.94 8.63 54.27 13.67 ;
      RECT  50.0 8.63 50.33 13.67 ;
      RECT  50.96 8.63 51.29 13.67 ;
      RECT  56.54 8.63 56.87 13.67 ;
      RECT  52.6 8.63 52.93 13.67 ;
      RECT  46.64 22.19 46.78 15.19 ;
      RECT  47.92 22.19 48.06 15.19 ;
      RECT  49.24 22.19 49.38 15.19 ;
      RECT  50.52 22.19 50.66 15.19 ;
      RECT  51.84 22.19 51.98 15.19 ;
      RECT  53.12 22.19 53.26 15.19 ;
      RECT  3.44 36.56 3.9 37.02 ;
      RECT  4.1 41.86 4.56 42.32 ;
      RECT  3.44 67.1 3.9 67.56 ;
      RECT  4.1 72.4 4.56 72.86 ;
      RECT  0.16 34.35 0.3 85.25 ;
      RECT  0.82 34.35 0.96 85.25 ;
      RECT  1.48 34.35 1.62 85.25 ;
      RECT  2.14 34.35 2.28 85.25 ;
      RECT  34.59 34.35 34.73 115.79 ;
      RECT  0.16 34.35 0.3 85.25 ;
      RECT  0.82 34.35 0.96 85.25 ;
      RECT  1.48 34.35 1.62 85.25 ;
      RECT  2.14 34.35 2.28 85.25 ;
      RECT  34.1 32.76 34.24 32.9 ;
      RECT  0.16 34.35 0.3 85.25 ;
      RECT  0.82 34.35 0.96 85.25 ;
      RECT  1.48 34.35 1.62 85.25 ;
      RECT  2.14 34.35 2.28 85.25 ;
      RECT  37.63 0.0 37.77 24.17 ;
      RECT  39.27 0.0 39.41 24.17 ;
      RECT  38.45 0.0 38.59 24.17 ;
      RECT  40.09 0.0 40.23 24.17 ;
      RECT  -55.0 -7.2 -54.66 -6.88 ;
      RECT  -46.1 -7.51 -45.78 -7.19 ;
      RECT  -55.78 -8.02 -55.47 -7.7 ;
      RECT  -55.0 -7.2 -54.66 -6.88 ;
      RECT  -33.53 -9.01 -33.39 -8.87 ;
      RECT  -37.3 -6.34 -37.16 -6.2 ;
      RECT  -55.78 -8.02 -55.47 -7.7 ;
      RECT  -55.0 -3.7 -54.66 -4.02 ;
      RECT  -46.1 -3.39 -45.78 -3.71 ;
      RECT  -55.78 -2.88 -55.47 -3.2 ;
      RECT  -55.0 -3.7 -54.66 -4.02 ;
      RECT  -33.53 -1.89 -33.39 -2.03 ;
      RECT  -37.3 -4.56 -37.16 -4.7 ;
      RECT  -55.78 -2.88 -55.47 -3.2 ;
      RECT  -55.0 -7.2 -54.66 -6.88 ;
      RECT  -55.0 -4.02 -54.66 -3.7 ;
      RECT  -33.53 -9.01 -33.39 -8.87 ;
      RECT  -37.3 -6.34 -37.16 -6.2 ;
      RECT  -33.53 -2.03 -33.39 -1.89 ;
      RECT  -37.3 -4.7 -37.16 -4.56 ;
      RECT  -55.78 -9.51 -55.64 -1.39 ;
      RECT  -40.68 24.17 -40.82 28.26 ;
      RECT  -53.75 24.17 -53.89 95.46 ;
      RECT  -55.0 -7.2 -54.66 -6.88 ;
      RECT  -55.0 -4.02 -54.66 -3.7 ;
      RECT  -25.11 -7.66 -24.97 -7.52 ;
      RECT  -40.82 24.17 -40.68 28.26 ;
      RECT  -19.57 20.98 -1.32 21.12 ;
      RECT  -17.28 8.54 -1.32 8.68 ;
      RECT  -17.44 12.86 -1.32 13.0 ;
      RECT  -12.59 4.75 -1.32 4.89 ;
      RECT  -7.18 -7.69 -1.32 -7.55 ;
      RECT  -12.8 103.28 -12.46 103.6 ;
      RECT  -3.9 102.97 -3.58 103.29 ;
      RECT  -13.58 102.46 -13.27 102.78 ;
      RECT  -12.8 106.78 -12.46 106.46 ;
      RECT  -3.9 107.09 -3.58 106.77 ;
      RECT  -13.58 107.6 -13.27 107.28 ;
      RECT  -12.8 111.4 -12.46 111.72 ;
      RECT  -3.9 111.09 -3.58 111.41 ;
      RECT  -13.58 110.58 -13.27 110.9 ;
      RECT  -12.8 114.9 -12.46 114.58 ;
      RECT  -3.9 115.21 -3.58 114.89 ;
      RECT  -13.58 115.72 -13.27 115.4 ;
      RECT  -12.8 103.28 -12.46 103.6 ;
      RECT  -12.8 106.46 -12.46 106.78 ;
      RECT  -12.8 111.4 -12.46 111.72 ;
      RECT  -12.8 114.58 -12.46 114.9 ;
      RECT  -3.9 102.97 -3.58 103.29 ;
      RECT  -3.9 106.77 -3.58 107.09 ;
      RECT  -3.9 111.09 -3.58 111.41 ;
      RECT  -3.9 114.89 -3.58 115.21 ;
      RECT  10.5 -7.2 10.84 -6.88 ;
      RECT  19.4 -7.51 19.72 -7.19 ;
      RECT  9.72 -8.02 10.03 -7.7 ;
      RECT  22.15 -7.2 22.49 -6.88 ;
      RECT  31.05 -7.51 31.37 -7.19 ;
      RECT  21.37 -8.02 21.68 -7.7 ;
      RECT  10.5 -7.2 10.84 -6.88 ;
      RECT  22.15 -7.2 22.49 -6.88 ;
      RECT  19.4 -7.51 19.72 -7.19 ;
      RECT  31.05 -7.51 31.37 -7.19 ;
   LAYER  m3 ;
      RECT  47.09 120.61 47.61 121.13 ;
      RECT  47.09 28.99 47.61 29.51 ;
      RECT  47.09 23.91 47.61 24.43 ;
      RECT  47.09 115.53 47.61 116.05 ;
      RECT  44.49 49.37 45.01 49.89 ;
      RECT  44.49 110.43 45.01 110.95 ;
      RECT  49.69 120.61 50.21 121.13 ;
      RECT  54.89 49.37 55.41 49.89 ;
      RECT  54.89 49.35 55.41 49.87 ;
      RECT  44.49 49.35 45.01 49.87 ;
      RECT  54.89 79.91 55.41 80.43 ;
      RECT  44.49 79.91 45.01 80.43 ;
      RECT  44.49 39.17 45.01 39.69 ;
      RECT  44.49 59.53 45.01 60.05 ;
      RECT  44.49 100.27 45.01 100.79 ;
      RECT  54.89 110.43 55.41 110.95 ;
      RECT  54.89 79.89 55.41 80.41 ;
      RECT  54.89 90.07 55.41 90.59 ;
      RECT  44.49 100.25 45.01 100.77 ;
      RECT  52.29 120.61 52.81 121.13 ;
      RECT  52.29 28.99 52.81 29.51 ;
      RECT  54.89 110.45 55.41 110.97 ;
      RECT  44.49 110.45 45.01 110.97 ;
      RECT  54.89 39.19 55.41 39.71 ;
      RECT  47.09 28.99 47.61 29.51 ;
      RECT  44.49 59.55 45.01 60.07 ;
      RECT  44.49 69.73 45.01 70.25 ;
      RECT  44.49 28.99 45.01 29.51 ;
      RECT  44.49 79.89 45.01 80.41 ;
      RECT  44.49 120.61 45.01 121.13 ;
      RECT  44.49 90.07 45.01 90.59 ;
      RECT  54.89 100.25 55.41 100.77 ;
      RECT  54.89 59.53 55.41 60.05 ;
      RECT  54.89 59.55 55.41 60.07 ;
      RECT  44.49 69.71 45.01 70.23 ;
      RECT  54.89 120.61 55.41 121.13 ;
      RECT  44.49 29.01 45.01 29.53 ;
      RECT  44.49 90.09 45.01 90.61 ;
      RECT  54.89 69.73 55.41 70.25 ;
      RECT  54.89 69.71 55.41 70.23 ;
      RECT  54.89 39.17 55.41 39.69 ;
      RECT  44.49 39.19 45.01 39.71 ;
      RECT  49.69 28.99 50.21 29.51 ;
      RECT  54.89 28.99 55.41 29.51 ;
      RECT  54.89 90.09 55.41 90.61 ;
      RECT  54.89 29.01 55.41 29.53 ;
      RECT  47.09 120.61 47.61 121.13 ;
      RECT  54.89 100.27 55.41 100.79 ;
      RECT  44.49 105.35 45.01 105.87 ;
      RECT  44.49 105.35 45.01 105.87 ;
      RECT  44.49 34.09 45.01 34.61 ;
      RECT  44.49 34.09 45.01 34.61 ;
      RECT  54.89 64.63 55.41 65.15 ;
      RECT  54.89 64.63 55.41 65.15 ;
      RECT  57.09 116.68 57.61 117.2 ;
      RECT  54.89 54.45 55.41 54.97 ;
      RECT  44.49 115.53 45.01 116.05 ;
      RECT  44.49 115.53 45.01 116.05 ;
      RECT  54.89 34.09 55.41 34.61 ;
      RECT  54.89 34.09 55.41 34.61 ;
      RECT  54.89 54.45 55.41 54.97 ;
      RECT  44.49 95.17 45.01 95.69 ;
      RECT  44.49 95.17 45.01 95.69 ;
      RECT  54.89 115.53 55.41 116.05 ;
      RECT  54.89 115.53 55.41 116.05 ;
      RECT  52.29 115.53 52.81 116.05 ;
      RECT  47.09 23.91 47.61 24.43 ;
      RECT  44.49 44.27 45.01 44.79 ;
      RECT  44.49 44.27 45.01 44.79 ;
      RECT  44.49 54.45 45.01 54.97 ;
      RECT  54.89 84.99 55.41 85.51 ;
      RECT  54.89 84.99 55.41 85.51 ;
      RECT  44.49 64.63 45.01 65.15 ;
      RECT  44.49 64.63 45.01 65.15 ;
      RECT  44.49 23.91 45.01 24.43 ;
      RECT  54.89 95.17 55.41 95.69 ;
      RECT  54.89 95.17 55.41 95.69 ;
      RECT  54.89 23.91 55.41 24.43 ;
      RECT  44.49 74.81 45.01 75.33 ;
      RECT  44.49 74.81 45.01 75.33 ;
      RECT  42.29 25.06 42.81 25.58 ;
      RECT  47.09 115.53 47.61 116.05 ;
      RECT  54.89 105.35 55.41 105.87 ;
      RECT  54.89 105.35 55.41 105.87 ;
      RECT  42.29 116.68 42.81 117.2 ;
      RECT  44.49 84.99 45.01 85.51 ;
      RECT  44.49 84.99 45.01 85.51 ;
      RECT  57.09 25.06 57.61 25.58 ;
      RECT  49.69 115.53 50.21 116.05 ;
      RECT  54.89 74.81 55.41 75.33 ;
      RECT  54.89 74.81 55.41 75.33 ;
      RECT  49.69 23.91 50.21 24.43 ;
      RECT  52.29 23.91 52.81 24.43 ;
      RECT  54.89 44.27 55.41 44.79 ;
      RECT  54.89 44.27 55.41 44.79 ;
      RECT  44.49 54.45 45.01 54.97 ;
      RECT  47.89 21.46 48.41 21.98 ;
      RECT  50.49 21.46 51.01 21.98 ;
      RECT  53.09 21.46 53.61 21.98 ;
      RECT  50.49 21.46 51.01 21.98 ;
      RECT  53.09 21.46 53.61 21.98 ;
      RECT  47.89 21.46 48.41 21.98 ;
      RECT  51.13 12.95 51.65 13.47 ;
      RECT  53.73 12.95 54.25 13.47 ;
      RECT  53.73 8.57 54.25 9.09 ;
      RECT  51.13 8.57 51.65 9.09 ;
      RECT  58.28 6.9 58.8 7.42 ;
      RECT  55.68 6.9 56.2 7.42 ;
      RECT  55.68 1.1 56.2 1.62 ;
      RECT  58.28 1.1 58.8 1.62 ;
      RECT  50.49 21.98 51.01 21.46 ;
      RECT  58.28 7.42 58.8 6.9 ;
      RECT  53.09 21.98 53.61 21.46 ;
      RECT  53.73 13.47 54.25 12.95 ;
      RECT  55.68 7.42 56.2 6.9 ;
      RECT  51.13 13.47 51.65 12.95 ;
      RECT  47.89 21.98 48.41 21.46 ;
      RECT  53.73 9.09 54.25 8.57 ;
      RECT  55.68 1.62 56.2 1.1 ;
      RECT  51.13 9.09 51.65 8.57 ;
      RECT  58.28 1.62 58.8 1.1 ;
      RECT  12.28 39.18 12.8 39.7 ;
      RECT  12.28 49.36 12.8 49.88 ;
      RECT  5.18 39.18 5.7 39.7 ;
      RECT  5.18 49.36 5.7 49.88 ;
      RECT  12.28 54.45 12.8 54.97 ;
      RECT  12.28 34.09 12.8 34.61 ;
      RECT  12.28 44.27 12.8 44.79 ;
      RECT  5.18 54.45 5.7 54.97 ;
      RECT  5.18 34.09 5.7 34.61 ;
      RECT  5.18 44.27 5.7 44.79 ;
      RECT  12.28 69.72 12.8 70.24 ;
      RECT  12.28 79.9 12.8 80.42 ;
      RECT  5.18 69.72 5.7 70.24 ;
      RECT  5.18 79.9 5.7 80.42 ;
      RECT  12.28 84.99 12.8 85.51 ;
      RECT  12.28 64.63 12.8 65.15 ;
      RECT  12.28 74.81 12.8 75.33 ;
      RECT  5.18 84.99 5.7 85.51 ;
      RECT  5.18 64.63 5.7 65.15 ;
      RECT  5.18 74.81 5.7 75.33 ;
      RECT  12.28 79.9 12.8 80.42 ;
      RECT  32.17 69.72 32.69 70.24 ;
      RECT  32.17 110.44 32.69 110.96 ;
      RECT  5.18 39.18 5.7 39.7 ;
      RECT  5.18 79.9 5.7 80.42 ;
      RECT  32.17 59.54 32.69 60.06 ;
      RECT  32.17 49.36 32.69 49.88 ;
      RECT  5.18 69.72 5.7 70.24 ;
      RECT  12.28 49.36 12.8 49.88 ;
      RECT  32.17 100.26 32.69 100.78 ;
      RECT  32.17 100.26 32.69 100.78 ;
      RECT  5.18 49.36 5.7 49.88 ;
      RECT  12.28 69.72 12.8 70.24 ;
      RECT  32.17 79.9 32.69 80.42 ;
      RECT  32.17 90.08 32.69 90.6 ;
      RECT  12.28 39.18 12.8 39.7 ;
      RECT  32.17 39.18 32.69 39.7 ;
      RECT  32.17 74.81 32.69 75.33 ;
      RECT  32.17 54.45 32.69 54.97 ;
      RECT  32.17 34.09 32.69 34.61 ;
      RECT  12.28 34.09 12.8 34.61 ;
      RECT  5.18 64.63 5.7 65.15 ;
      RECT  5.18 34.09 5.7 34.61 ;
      RECT  12.28 54.45 12.8 54.97 ;
      RECT  12.28 64.63 12.8 65.15 ;
      RECT  32.17 95.17 32.69 95.69 ;
      RECT  5.18 54.45 5.7 54.97 ;
      RECT  12.28 44.27 12.8 44.79 ;
      RECT  32.17 115.53 32.69 116.05 ;
      RECT  32.17 84.99 32.69 85.51 ;
      RECT  12.28 84.99 12.8 85.51 ;
      RECT  5.18 74.81 5.7 75.33 ;
      RECT  5.18 44.27 5.7 44.79 ;
      RECT  32.17 105.35 32.69 105.87 ;
      RECT  32.17 44.27 32.69 44.79 ;
      RECT  12.28 74.81 12.8 75.33 ;
      RECT  32.17 64.63 32.69 65.15 ;
      RECT  5.18 84.99 5.7 85.51 ;
      RECT  39.04 59.54 39.56 60.06 ;
      RECT  39.04 79.9 39.56 80.42 ;
      RECT  39.04 39.18 39.56 39.7 ;
      RECT  39.04 69.72 39.56 70.24 ;
      RECT  39.04 90.08 39.56 90.6 ;
      RECT  39.04 110.44 39.56 110.96 ;
      RECT  39.04 100.26 39.56 100.78 ;
      RECT  39.04 100.26 39.56 100.78 ;
      RECT  39.04 49.36 39.56 49.88 ;
      RECT  39.04 54.45 39.56 54.97 ;
      RECT  39.04 44.27 39.56 44.79 ;
      RECT  39.04 74.81 39.56 75.33 ;
      RECT  39.04 95.17 39.56 95.69 ;
      RECT  39.04 34.09 39.56 34.61 ;
      RECT  39.04 115.53 39.56 116.05 ;
      RECT  39.04 84.99 39.56 85.51 ;
      RECT  39.04 105.35 39.56 105.87 ;
      RECT  39.04 64.63 39.56 65.15 ;
      RECT  39.04 90.08 39.56 90.6 ;
      RECT  32.17 29.0 32.69 29.52 ;
      RECT  39.04 59.54 39.56 60.06 ;
      RECT  39.04 69.72 39.56 70.24 ;
      RECT  12.28 39.18 12.8 39.7 ;
      RECT  12.28 49.36 12.8 49.88 ;
      RECT  39.04 39.18 39.56 39.7 ;
      RECT  39.04 110.44 39.56 110.96 ;
      RECT  5.18 39.18 5.7 39.7 ;
      RECT  5.18 49.36 5.7 49.88 ;
      RECT  5.18 79.9 5.7 80.42 ;
      RECT  32.17 100.26 32.69 100.78 ;
      RECT  5.18 69.72 5.7 70.24 ;
      RECT  39.04 49.36 39.56 49.88 ;
      RECT  32.17 69.72 32.69 70.24 ;
      RECT  32.17 90.08 32.69 90.6 ;
      RECT  32.17 39.18 32.69 39.7 ;
      RECT  12.28 79.9 12.8 80.42 ;
      RECT  32.7 30.93 33.22 31.45 ;
      RECT  32.17 110.44 32.69 110.96 ;
      RECT  32.17 79.9 32.69 80.42 ;
      RECT  39.04 100.26 39.56 100.78 ;
      RECT  32.17 49.36 32.69 49.88 ;
      RECT  39.04 79.9 39.56 80.42 ;
      RECT  32.17 59.54 32.69 60.06 ;
      RECT  12.28 69.72 12.8 70.24 ;
      RECT  5.18 64.63 5.7 65.15 ;
      RECT  5.18 44.27 5.7 44.79 ;
      RECT  32.17 74.81 32.69 75.33 ;
      RECT  32.17 34.09 32.69 34.61 ;
      RECT  32.17 54.45 32.69 54.97 ;
      RECT  39.04 64.63 39.56 65.15 ;
      RECT  12.28 34.09 12.8 34.61 ;
      RECT  39.04 84.99 39.56 85.51 ;
      RECT  32.17 64.63 32.69 65.15 ;
      RECT  32.17 115.53 32.69 116.05 ;
      RECT  5.18 54.45 5.7 54.97 ;
      RECT  39.04 105.35 39.56 105.87 ;
      RECT  32.17 105.35 32.69 105.87 ;
      RECT  12.28 54.45 12.8 54.97 ;
      RECT  12.28 84.99 12.8 85.51 ;
      RECT  12.28 44.27 12.8 44.79 ;
      RECT  39.04 115.53 39.56 116.05 ;
      RECT  12.28 74.81 12.8 75.33 ;
      RECT  39.04 34.09 39.56 34.61 ;
      RECT  5.18 74.81 5.7 75.33 ;
      RECT  39.04 74.81 39.56 75.33 ;
      RECT  5.18 34.09 5.7 34.61 ;
      RECT  5.18 84.99 5.7 85.51 ;
      RECT  39.04 54.45 39.56 54.97 ;
      RECT  32.17 95.17 32.69 95.69 ;
      RECT  12.28 64.63 12.8 65.15 ;
      RECT  32.17 84.99 32.69 85.51 ;
      RECT  32.17 44.27 32.69 44.79 ;
      RECT  39.04 44.27 39.56 44.79 ;
      RECT  39.04 95.17 39.56 95.69 ;
      RECT  0.0 14.22 46.71 14.52 ;
      RECT  50.49 21.46 51.01 21.98 ;
      RECT  44.49 49.37 45.01 49.89 ;
      RECT  12.28 49.36 12.8 49.88 ;
      RECT  49.69 120.61 50.21 121.13 ;
      RECT  44.49 79.91 45.01 80.43 ;
      RECT  53.09 21.46 53.61 21.98 ;
      RECT  51.13 12.95 51.65 13.47 ;
      RECT  39.04 79.9 39.56 80.42 ;
      RECT  52.29 120.61 52.81 121.13 ;
      RECT  32.17 110.44 32.69 110.96 ;
      RECT  52.29 28.99 52.81 29.51 ;
      RECT  44.49 59.55 45.01 60.07 ;
      RECT  44.49 90.07 45.01 90.59 ;
      RECT  44.49 69.71 45.01 70.23 ;
      RECT  54.89 69.73 55.41 70.25 ;
      RECT  44.49 39.19 45.01 39.71 ;
      RECT  54.89 100.27 55.41 100.79 ;
      RECT  54.89 49.37 55.41 49.89 ;
      RECT  44.49 49.35 45.01 49.87 ;
      RECT  54.89 79.91 55.41 80.43 ;
      RECT  32.7 30.93 33.22 31.45 ;
      RECT  32.17 69.72 32.69 70.24 ;
      RECT  58.28 6.9 58.8 7.42 ;
      RECT  54.89 90.07 55.41 90.59 ;
      RECT  54.89 79.89 55.41 80.41 ;
      RECT  39.04 110.44 39.56 110.96 ;
      RECT  44.49 69.73 45.01 70.25 ;
      RECT  44.49 28.99 45.01 29.51 ;
      RECT  54.89 59.53 55.41 60.05 ;
      RECT  54.89 59.55 55.41 60.07 ;
      RECT  39.04 59.54 39.56 60.06 ;
      RECT  54.89 69.71 55.41 70.23 ;
      RECT  44.49 90.09 45.01 90.61 ;
      RECT  49.69 28.99 50.21 29.51 ;
      RECT  54.89 90.09 55.41 90.61 ;
      RECT  39.04 100.26 39.56 100.78 ;
      RECT  12.28 69.72 12.8 70.24 ;
      RECT  12.28 39.18 12.8 39.7 ;
      RECT  54.89 49.35 55.41 49.87 ;
      RECT  5.18 49.36 5.7 49.88 ;
      RECT  5.18 79.9 5.7 80.42 ;
      RECT  54.89 100.25 55.41 100.77 ;
      RECT  55.68 6.9 56.2 7.42 ;
      RECT  39.04 90.08 39.56 90.6 ;
      RECT  32.17 100.26 32.69 100.78 ;
      RECT  5.18 69.72 5.7 70.24 ;
      RECT  32.17 59.54 32.69 60.06 ;
      RECT  44.49 29.01 45.01 29.53 ;
      RECT  54.89 28.99 55.41 29.51 ;
      RECT  47.89 21.46 48.41 21.98 ;
      RECT  44.49 110.43 45.01 110.95 ;
      RECT  32.17 39.18 32.69 39.7 ;
      RECT  39.04 49.36 39.56 49.88 ;
      RECT  32.17 29.0 32.69 29.52 ;
      RECT  44.49 39.17 45.01 39.69 ;
      RECT  44.49 59.53 45.01 60.05 ;
      RECT  39.04 69.72 39.56 70.24 ;
      RECT  5.18 39.18 5.7 39.7 ;
      RECT  32.17 49.36 32.69 49.88 ;
      RECT  44.49 100.27 45.01 100.79 ;
      RECT  54.89 110.43 55.41 110.95 ;
      RECT  44.49 100.25 45.01 100.77 ;
      RECT  32.17 79.9 32.69 80.42 ;
      RECT  12.28 79.9 12.8 80.42 ;
      RECT  44.49 110.45 45.01 110.97 ;
      RECT  54.89 39.19 55.41 39.71 ;
      RECT  47.09 28.99 47.61 29.51 ;
      RECT  44.49 79.89 45.01 80.41 ;
      RECT  44.49 120.61 45.01 121.13 ;
      RECT  32.17 90.08 32.69 90.6 ;
      RECT  39.04 39.18 39.56 39.7 ;
      RECT  53.73 12.95 54.25 13.47 ;
      RECT  54.89 120.61 55.41 121.13 ;
      RECT  54.89 39.17 55.41 39.69 ;
      RECT  54.89 110.45 55.41 110.97 ;
      RECT  54.89 29.01 55.41 29.53 ;
      RECT  47.09 120.61 47.61 121.13 ;
      RECT  44.49 105.35 45.01 105.87 ;
      RECT  39.04 54.45 39.56 54.97 ;
      RECT  44.49 34.09 45.01 34.61 ;
      RECT  39.04 64.63 39.56 65.15 ;
      RECT  32.17 64.63 32.69 65.15 ;
      RECT  39.04 115.53 39.56 116.05 ;
      RECT  32.17 84.99 32.69 85.51 ;
      RECT  5.18 44.27 5.7 44.79 ;
      RECT  5.18 84.99 5.7 85.51 ;
      RECT  12.28 54.45 12.8 54.97 ;
      RECT  54.89 64.63 55.41 65.15 ;
      RECT  57.09 116.68 57.61 117.2 ;
      RECT  54.89 54.45 55.41 54.97 ;
      RECT  44.49 115.53 45.01 116.05 ;
      RECT  32.17 115.53 32.69 116.05 ;
      RECT  54.89 34.09 55.41 34.61 ;
      RECT  44.49 95.17 45.01 95.69 ;
      RECT  54.89 115.53 55.41 116.05 ;
      RECT  52.29 115.53 52.81 116.05 ;
      RECT  47.09 23.91 47.61 24.43 ;
      RECT  53.73 8.57 54.25 9.09 ;
      RECT  44.49 44.27 45.01 44.79 ;
      RECT  5.18 54.45 5.7 54.97 ;
      RECT  12.28 64.63 12.8 65.15 ;
      RECT  32.17 105.35 32.69 105.87 ;
      RECT  54.89 84.99 55.41 85.51 ;
      RECT  32.17 95.17 32.69 95.69 ;
      RECT  39.04 95.17 39.56 95.69 ;
      RECT  44.49 64.63 45.01 65.15 ;
      RECT  32.17 34.09 32.69 34.61 ;
      RECT  54.89 95.17 55.41 95.69 ;
      RECT  44.49 23.91 45.01 24.43 ;
      RECT  51.13 8.57 51.65 9.09 ;
      RECT  54.89 23.91 55.41 24.43 ;
      RECT  12.28 44.27 12.8 44.79 ;
      RECT  32.17 44.27 32.69 44.79 ;
      RECT  44.49 74.81 45.01 75.33 ;
      RECT  58.28 1.1 58.8 1.62 ;
      RECT  42.29 25.06 42.81 25.58 ;
      RECT  5.18 34.09 5.7 34.61 ;
      RECT  47.09 115.53 47.61 116.05 ;
      RECT  55.68 1.1 56.2 1.62 ;
      RECT  39.04 84.99 39.56 85.51 ;
      RECT  39.04 74.81 39.56 75.33 ;
      RECT  54.89 105.35 55.41 105.87 ;
      RECT  42.29 116.68 42.81 117.2 ;
      RECT  5.18 64.63 5.7 65.15 ;
      RECT  44.49 84.99 45.01 85.51 ;
      RECT  32.17 54.45 32.69 54.97 ;
      RECT  32.17 74.81 32.69 75.33 ;
      RECT  57.09 25.06 57.61 25.58 ;
      RECT  49.69 115.53 50.21 116.05 ;
      RECT  5.18 74.81 5.7 75.33 ;
      RECT  54.89 74.81 55.41 75.33 ;
      RECT  12.28 34.09 12.8 34.61 ;
      RECT  49.69 23.91 50.21 24.43 ;
      RECT  52.29 23.91 52.81 24.43 ;
      RECT  54.89 44.27 55.41 44.79 ;
      RECT  39.04 34.09 39.56 34.61 ;
      RECT  39.04 44.27 39.56 44.79 ;
      RECT  39.04 105.35 39.56 105.87 ;
      RECT  12.28 74.81 12.8 75.33 ;
      RECT  12.28 84.99 12.8 85.51 ;
      RECT  44.49 54.45 45.01 54.97 ;
      RECT  -56.49 -5.71 -55.97 -5.19 ;
      RECT  -56.49 -5.71 -55.97 -5.19 ;
      RECT  -56.49 -1.63 -55.97 -1.11 ;
      RECT  -56.49 -9.79 -55.97 -9.27 ;
      RECT  -51.17 32.31 -51.69 32.83 ;
      RECT  -51.17 65.91 -51.69 66.43 ;
      RECT  -51.17 99.51 -51.69 100.03 ;
      RECT  -44.89 32.31 -45.41 32.83 ;
      RECT  -44.89 99.51 -45.41 100.03 ;
      RECT  -51.17 82.71 -51.69 83.23 ;
      RECT  -44.89 49.11 -45.41 49.63 ;
      RECT  -44.89 82.71 -45.41 83.23 ;
      RECT  -44.89 65.91 -45.41 66.43 ;
      RECT  -51.17 49.11 -51.69 49.63 ;
      RECT  -44.89 23.91 -45.41 24.43 ;
      RECT  -51.17 57.51 -51.69 58.03 ;
      RECT  -51.17 40.71 -51.69 41.23 ;
      RECT  -51.17 23.91 -51.69 24.43 ;
      RECT  -51.17 91.11 -51.69 91.63 ;
      RECT  -44.89 40.71 -45.41 41.23 ;
      RECT  -44.89 74.31 -45.41 74.83 ;
      RECT  -44.89 57.51 -45.41 58.03 ;
      RECT  -44.89 91.11 -45.41 91.63 ;
      RECT  -51.17 74.31 -51.69 74.83 ;
      RECT  -51.69 99.51 -51.17 100.03 ;
      RECT  -45.41 82.71 -44.89 83.23 ;
      RECT  -45.41 65.91 -44.89 66.43 ;
      RECT  -45.41 99.51 -44.89 100.03 ;
      RECT  -51.69 49.11 -51.17 49.63 ;
      RECT  -51.69 65.91 -51.17 66.43 ;
      RECT  -45.41 32.31 -44.89 32.83 ;
      RECT  -45.41 49.11 -44.89 49.63 ;
      RECT  -56.49 -5.71 -55.97 -5.19 ;
      RECT  -51.69 82.71 -51.17 83.23 ;
      RECT  -51.69 32.31 -51.17 32.83 ;
      RECT  -51.69 57.51 -51.17 58.03 ;
      RECT  -51.69 23.91 -51.17 24.43 ;
      RECT  -45.41 74.31 -44.89 74.83 ;
      RECT  -45.41 57.51 -44.89 58.03 ;
      RECT  -56.49 -1.63 -55.97 -1.11 ;
      RECT  -45.41 40.71 -44.89 41.23 ;
      RECT  -51.69 91.11 -51.17 91.63 ;
      RECT  -51.69 40.71 -51.17 41.23 ;
      RECT  -45.41 91.11 -44.89 91.63 ;
      RECT  -45.41 23.91 -44.89 24.43 ;
      RECT  -51.69 74.31 -51.17 74.83 ;
      RECT  -56.49 -9.79 -55.97 -9.27 ;
      RECT  -12.97 102.76 -1.32 103.06 ;
      RECT  -7.93 112.89 -7.41 113.41 ;
      RECT  -7.93 104.77 -7.41 105.29 ;
      RECT  -7.93 104.77 -7.41 105.29 ;
      RECT  -7.93 112.89 -7.41 113.41 ;
      RECT  -7.93 108.81 -7.41 109.33 ;
      RECT  -7.93 116.97 -7.41 117.49 ;
      RECT  -7.93 100.69 -7.41 101.21 ;
      RECT  -7.93 108.85 -7.41 109.37 ;
      RECT  10.33 -7.72 33.63 -7.42 ;
      RECT  27.01 -5.71 27.53 -5.19 ;
      RECT  15.37 -5.71 15.89 -5.19 ;
      RECT  27.01 -9.79 27.53 -9.27 ;
      RECT  15.37 -9.79 15.89 -9.27 ;
   LAYER  m4 ;
   END
   END    sram_2_16_sky130A
END    LIBRARY
