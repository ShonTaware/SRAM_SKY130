SRAM Cell N Curve

.lib "./libs/models/sky130.lib.spice" tt

*** Inverter 1
XM1 qbar q gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.21
XM2 qbar q vdd vdd sky130_fd_pr__pfet_01v8 w=0.84 l=0.21

*** Inverter 2 
XM3 q qbar gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.21
XM4 q qbar vdd vdd sky130_fd_pr__pfet_01v8 w=0.84 l=0.21


*** Access Transistors
XM5 bl wl q gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.21
XM6 blbar wl qbar gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.21

V1 vdd gnd dc 1.8V
Vin Q gnd dc 1.8V
Vwl wl gnd dc 1.8v
Vbl bl gnd dc 1.8v
Vblbar blbar gnd dc 1.8v

.dc Vin 0 1.8 0.01
.control
run
plot -I(Vin)
.endc
.end

