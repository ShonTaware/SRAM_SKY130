magic
tech sky130A
timestamp 1613393172
<< fence >>
rect 1 -240 586 178
<< nwell >>
rect 1 -19 481 178
<< nmos >>
rect 68 -135 83 -93
rect 232 -135 247 -93
rect 372 -132 387 -77
rect 517 -93 559 -78
<< pmos >>
rect 68 15 83 57
rect 232 15 247 57
rect 372 2 387 57
<< ndiff >>
rect 330 -93 372 -77
rect 25 -114 68 -93
rect 25 -131 32 -114
rect 49 -131 68 -114
rect 25 -135 68 -131
rect 83 -97 126 -93
rect 83 -114 100 -97
rect 117 -114 126 -97
rect 83 -135 126 -114
rect 189 -114 232 -93
rect 189 -131 197 -114
rect 214 -131 232 -114
rect 189 -135 232 -131
rect 247 -97 290 -93
rect 247 -114 265 -97
rect 282 -114 290 -97
rect 247 -135 290 -114
rect 330 -110 339 -93
rect 356 -110 372 -93
rect 330 -132 372 -110
rect 387 -93 431 -77
rect 517 -40 559 -36
rect 517 -57 528 -40
rect 545 -57 559 -40
rect 517 -78 559 -57
rect 387 -110 404 -93
rect 421 -110 431 -93
rect 387 -132 431 -110
rect 517 -115 559 -93
rect 517 -132 531 -115
rect 548 -132 559 -115
rect 517 -137 559 -132
<< pdiff >>
rect 25 42 68 57
rect 25 25 32 42
rect 49 25 68 42
rect 25 15 68 25
rect 83 45 126 57
rect 83 28 99 45
rect 116 28 126 45
rect 83 15 126 28
rect 189 43 232 57
rect 189 26 197 43
rect 214 26 232 43
rect 189 15 232 26
rect 247 43 290 57
rect 247 26 263 43
rect 280 26 290 43
rect 247 15 290 26
rect 330 30 372 57
rect 330 13 338 30
rect 355 13 372 30
rect 330 2 372 13
rect 387 44 431 57
rect 387 30 432 44
rect 387 13 409 30
rect 426 13 432 30
rect 387 2 432 13
<< ndiffc >>
rect 32 -131 49 -114
rect 100 -114 117 -97
rect 197 -131 214 -114
rect 265 -114 282 -97
rect 339 -110 356 -93
rect 528 -57 545 -40
rect 404 -110 421 -93
rect 531 -132 548 -115
<< pdiffc >>
rect 32 25 49 42
rect 99 28 116 45
rect 197 26 214 43
rect 263 26 280 43
rect 338 13 355 30
rect 409 13 426 30
<< psubdiff >>
rect 24 -234 58 -217
rect 75 -234 93 -217
rect 141 -234 165 -217
rect 182 -234 221 -217
rect 480 -233 496 -216
rect 513 -233 560 -216
<< nsubdiff >>
rect 25 141 66 158
rect 83 141 98 158
rect 159 141 172 158
rect 189 141 223 158
<< psubdiffcont >>
rect 58 -234 75 -217
rect 165 -234 182 -217
rect 496 -233 513 -216
<< nsubdiffcont >>
rect 66 141 83 158
rect 172 141 189 158
<< poly >>
rect 362 98 397 104
rect 362 81 372 98
rect 389 81 397 98
rect 68 57 83 70
rect 232 57 247 70
rect 362 69 397 81
rect 372 57 387 69
rect 68 -29 83 15
rect 232 -26 247 15
rect 372 -8 387 2
rect 372 -23 504 -8
rect 38 -37 83 -29
rect 38 -54 46 -37
rect 63 -54 83 -37
rect 38 -62 83 -54
rect 202 -34 247 -26
rect 202 -51 209 -34
rect 226 -51 247 -34
rect 202 -59 247 -51
rect 68 -93 83 -62
rect 232 -93 247 -59
rect 372 -77 387 -63
rect 489 -78 504 -23
rect 489 -93 517 -78
rect 559 -93 572 -78
rect 68 -148 83 -135
rect 232 -148 247 -135
rect 372 -145 387 -132
rect 362 -153 397 -145
rect 362 -170 371 -153
rect 388 -170 397 -153
rect 362 -180 397 -170
<< polycont >>
rect 372 81 389 98
rect 46 -54 63 -37
rect 209 -51 226 -34
rect 371 -170 388 -153
<< locali >>
rect 25 141 33 158
rect 50 141 66 158
rect 83 141 98 158
rect 159 141 172 158
rect 189 141 195 158
rect 212 141 223 158
rect 33 57 50 141
rect 195 57 212 141
rect 362 98 397 104
rect 362 81 372 98
rect 389 81 397 98
rect 362 69 397 81
rect 25 42 60 57
rect 25 25 32 42
rect 49 25 60 42
rect 25 15 60 25
rect 91 45 126 57
rect 91 28 99 45
rect 116 28 126 45
rect 91 15 126 28
rect 189 43 224 57
rect 189 26 197 43
rect 214 26 224 43
rect 189 15 224 26
rect 255 43 290 57
rect 255 26 263 43
rect 280 26 290 43
rect 255 15 290 26
rect 330 30 365 44
rect 109 7 126 15
rect 266 7 283 15
rect 330 13 338 30
rect 355 13 365 30
rect 330 2 365 13
rect 397 30 432 44
rect 397 13 409 30
rect 426 13 432 30
rect 397 2 432 13
rect 38 -37 68 -29
rect 19 -54 46 -37
rect 63 -54 68 -37
rect 38 -62 68 -54
rect 202 -34 232 -26
rect 202 -51 209 -34
rect 226 -51 232 -34
rect 202 -59 232 -51
rect 340 -36 357 2
rect 109 -93 126 -87
rect 340 -77 357 -53
rect 409 -36 426 2
rect 409 -40 586 -36
rect 409 -53 528 -40
rect 409 -77 426 -53
rect 517 -57 528 -53
rect 545 -53 586 -40
rect 545 -57 559 -53
rect 517 -61 559 -57
rect 266 -93 283 -86
rect 330 -93 365 -77
rect 91 -97 126 -93
rect 25 -114 60 -106
rect 25 -131 32 -114
rect 49 -131 60 -114
rect 91 -114 100 -97
rect 117 -114 126 -97
rect 255 -97 290 -93
rect 91 -118 126 -114
rect 189 -114 224 -110
rect 25 -135 60 -131
rect 189 -131 197 -114
rect 214 -131 224 -114
rect 255 -114 265 -97
rect 282 -114 290 -97
rect 255 -118 290 -114
rect 330 -110 339 -93
rect 356 -110 365 -93
rect 330 -119 365 -110
rect 396 -93 431 -77
rect 396 -110 404 -93
rect 421 -110 431 -93
rect 396 -119 431 -110
rect 517 -115 559 -112
rect 189 -135 224 -131
rect 517 -132 531 -115
rect 548 -132 559 -115
rect 32 -217 49 -135
rect 197 -217 214 -135
rect 517 -137 559 -132
rect 362 -153 397 -145
rect 362 -170 371 -153
rect 388 -170 397 -153
rect 362 -180 397 -170
rect 525 -216 542 -137
rect 24 -234 32 -217
rect 49 -234 58 -217
rect 75 -234 93 -217
rect 141 -234 165 -217
rect 182 -234 197 -217
rect 214 -234 221 -217
rect 480 -233 496 -216
rect 513 -233 525 -216
rect 542 -233 560 -216
<< viali >>
rect 33 141 50 158
rect 195 141 212 158
rect 372 81 389 98
rect 109 -10 126 7
rect 266 -10 283 7
rect 209 -51 226 -34
rect 340 -53 357 -36
rect 109 -87 126 -69
rect 266 -86 283 -69
rect 371 -170 388 -153
rect 32 -234 49 -217
rect 197 -234 214 -217
rect 525 -233 542 -216
<< metal1 >>
rect 22 158 223 164
rect 22 141 33 158
rect 50 141 195 158
rect 212 141 223 158
rect 22 135 223 141
rect 362 98 397 120
rect 362 81 372 98
rect 389 81 397 98
rect 362 69 397 81
rect 103 7 132 14
rect 103 -10 109 7
rect 126 -10 132 7
rect 103 -25 132 -10
rect 260 7 289 13
rect 260 -10 266 7
rect 283 -10 289 7
rect 103 -34 231 -25
rect 103 -51 209 -34
rect 226 -51 231 -34
rect 103 -59 231 -51
rect 260 -30 289 -10
rect 260 -36 364 -30
rect 260 -53 340 -36
rect 357 -53 364 -36
rect 260 -59 364 -53
rect 103 -69 132 -59
rect 103 -87 109 -69
rect 126 -87 132 -69
rect 103 -93 132 -87
rect 260 -69 289 -59
rect 260 -86 266 -69
rect 283 -86 289 -69
rect 260 -92 289 -86
rect 359 -153 416 -147
rect 359 -170 371 -153
rect 388 -170 416 -153
rect 359 -176 416 -170
rect 22 -216 567 -211
rect 22 -217 525 -216
rect 22 -234 32 -217
rect 49 -234 197 -217
rect 214 -233 525 -217
rect 542 -233 567 -216
rect 214 -234 567 -233
rect 22 -240 567 -234
<< labels >>
flabel locali 19 -53 37 -38 0 FreeSans 152 0 0 0 in
flabel locali 424 -52 458 -37 0 FreeSans 152 0 0 0 out
flabel metal1 82 -233 125 -218 0 FreeSans 152 0 0 0 gnd
flabel metal1 146 -49 163 -32 0 FreeSans 120 0 0 0 inb
flabel metal1 294 -51 316 -38 0 FreeSans 120 0 0 0 out1
flabel metal1 109 141 137 157 0 FreeSans 152 0 0 0 vdd
flabel metal1 399 -169 416 -152 0 FreeSans 120 0 0 0 en
flabel metal1 371 109 387 118 0 FreeSans 120 0 0 0 enb
<< end >>
