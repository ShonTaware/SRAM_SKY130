magic
tech sky130A
timestamp 1615997386
<< nwell >>
rect -106 271 1165 451
<< nmos >>
rect -42 55 -27 97
rect 101 55 116 97
rect 222 55 237 97
rect 393 55 408 97
rect 488 55 503 97
rect 681 55 696 97
rect 802 55 817 97
rect 997 55 1012 97
rect 1092 55 1107 97
<< pmos >>
rect -42 289 -27 344
rect 101 289 116 344
rect 222 289 237 344
rect 393 289 408 344
rect 488 289 503 344
rect 681 289 696 344
rect 802 289 817 344
rect 997 289 1012 344
rect 1092 289 1107 344
<< ndiff >>
rect -88 86 -42 97
rect -88 69 -78 86
rect -61 69 -42 86
rect -88 55 -42 69
rect -27 86 19 97
rect -27 69 -9 86
rect 8 69 19 86
rect -27 55 19 69
rect 55 86 101 97
rect 55 69 65 86
rect 82 69 101 86
rect 55 55 101 69
rect 116 86 222 97
rect 116 69 175 86
rect 192 69 222 86
rect 116 55 222 69
rect 237 86 305 97
rect 237 69 270 86
rect 287 69 305 86
rect 237 55 305 69
rect 340 85 393 97
rect 340 68 353 85
rect 370 68 393 85
rect 340 55 393 68
rect 408 86 488 97
rect 408 69 441 86
rect 458 69 488 86
rect 408 55 488 69
rect 503 86 565 97
rect 503 69 516 86
rect 533 69 565 86
rect 503 55 565 69
rect 616 86 681 97
rect 616 69 645 86
rect 662 69 681 86
rect 616 55 681 69
rect 696 86 802 97
rect 696 69 755 86
rect 772 69 802 86
rect 696 55 802 69
rect 817 86 896 97
rect 817 69 850 86
rect 867 69 896 86
rect 817 55 896 69
rect 941 86 997 97
rect 941 69 957 86
rect 974 69 997 86
rect 941 55 997 69
rect 1012 86 1092 97
rect 1012 69 1045 86
rect 1062 69 1092 86
rect 1012 55 1092 69
rect 1107 86 1147 97
rect 1107 69 1120 86
rect 1137 69 1147 86
rect 1107 55 1147 69
<< pdiff >>
rect -88 326 -42 344
rect -88 309 -78 326
rect -61 309 -42 326
rect -88 289 -42 309
rect -27 326 19 344
rect -27 309 -9 326
rect 8 309 19 326
rect -27 289 19 309
rect 55 326 101 344
rect 55 309 65 326
rect 82 309 101 326
rect 55 289 101 309
rect 116 326 222 344
rect 116 309 175 326
rect 192 309 222 326
rect 116 289 222 309
rect 237 326 305 344
rect 237 309 270 326
rect 287 309 305 326
rect 237 289 305 309
rect 340 326 393 344
rect 340 309 358 326
rect 375 309 393 326
rect 340 289 393 309
rect 408 326 488 344
rect 408 309 441 326
rect 458 309 488 326
rect 408 289 488 309
rect 503 326 566 344
rect 503 309 516 326
rect 533 309 566 326
rect 503 289 566 309
rect 617 326 681 344
rect 617 309 645 326
rect 662 309 681 326
rect 617 289 681 309
rect 696 326 802 344
rect 696 309 755 326
rect 772 309 802 326
rect 696 289 802 309
rect 817 326 896 344
rect 817 309 850 326
rect 867 309 896 326
rect 817 289 896 309
rect 941 326 997 344
rect 941 309 954 326
rect 971 309 997 326
rect 941 289 997 309
rect 1012 326 1092 344
rect 1012 309 1045 326
rect 1062 309 1092 326
rect 1012 289 1092 309
rect 1107 326 1147 344
rect 1107 309 1120 326
rect 1137 309 1147 326
rect 1107 289 1147 309
<< ndiffc >>
rect -78 69 -61 86
rect -9 69 8 86
rect 65 69 82 86
rect 175 69 192 86
rect 270 69 287 86
rect 353 68 370 85
rect 441 69 458 86
rect 516 69 533 86
rect 645 69 662 86
rect 755 69 772 86
rect 850 69 867 86
rect 957 69 974 86
rect 1045 69 1062 86
rect 1120 69 1137 86
<< pdiffc >>
rect -78 309 -61 326
rect -9 309 8 326
rect 65 309 82 326
rect 175 309 192 326
rect 270 309 287 326
rect 358 309 375 326
rect 441 309 458 326
rect 516 309 533 326
rect 645 309 662 326
rect 755 309 772 326
rect 850 309 867 326
rect 954 309 971 326
rect 1045 309 1062 326
rect 1120 309 1137 326
<< psubdiff >>
rect -103 6 -62 18
rect -103 -11 -91 6
rect -74 -11 -62 6
rect -103 -23 -62 -11
rect 40 6 81 18
rect 40 -11 52 6
rect 69 -11 81 6
rect 40 -23 81 -11
rect 144 6 185 18
rect 144 -11 156 6
rect 173 -11 185 6
rect 144 -23 185 -11
rect 255 6 296 18
rect 255 -11 267 6
rect 284 -11 296 6
rect 255 -23 296 -11
rect 440 6 481 18
rect 440 -11 452 6
rect 469 -11 481 6
rect 440 -23 481 -11
rect 620 6 661 18
rect 620 -11 632 6
rect 649 -11 661 6
rect 620 -23 661 -11
rect 724 6 765 18
rect 724 -11 736 6
rect 753 -11 765 6
rect 724 -23 765 -11
rect 835 6 876 18
rect 835 -11 847 6
rect 864 -11 876 6
rect 835 -23 876 -11
rect 1044 6 1085 18
rect 1044 -11 1056 6
rect 1073 -11 1085 6
rect 1044 -23 1085 -11
<< nsubdiff >>
rect -88 415 -35 433
rect -88 398 -70 415
rect -53 398 -35 415
rect -88 380 -35 398
rect 55 415 108 433
rect 55 398 73 415
rect 90 398 108 415
rect 55 380 108 398
rect 207 415 260 433
rect 207 398 225 415
rect 242 398 260 415
rect 207 380 260 398
rect 441 415 494 433
rect 441 398 459 415
rect 476 398 494 415
rect 441 380 494 398
rect 635 415 688 433
rect 635 398 653 415
rect 670 398 688 415
rect 635 380 688 398
rect 787 415 840 433
rect 787 398 805 415
rect 822 398 840 415
rect 787 380 840 398
rect 1045 415 1098 433
rect 1045 398 1063 415
rect 1080 398 1098 415
rect 1045 380 1098 398
<< psubdiffcont >>
rect -91 -11 -74 6
rect 52 -11 69 6
rect 156 -11 173 6
rect 267 -11 284 6
rect 452 -11 469 6
rect 632 -11 649 6
rect 736 -11 753 6
rect 847 -11 864 6
rect 1056 -11 1073 6
<< nsubdiffcont >>
rect -70 398 -53 415
rect 73 398 90 415
rect 225 398 242 415
rect 459 398 476 415
rect 653 398 670 415
rect 805 398 822 415
rect 1063 398 1080 415
<< poly >>
rect -42 344 -27 359
rect 101 344 116 359
rect 222 344 237 359
rect 393 344 408 359
rect 488 344 503 359
rect 681 344 696 359
rect 802 344 817 359
rect 997 344 1012 359
rect 1092 344 1107 359
rect -98 216 -65 224
rect -98 199 -90 216
rect -73 215 -65 216
rect -42 217 -27 289
rect 101 217 116 289
rect 222 267 237 289
rect 393 269 408 289
rect 213 259 246 267
rect 213 242 221 259
rect 238 242 246 259
rect 213 234 246 242
rect 393 261 426 269
rect 393 244 401 261
rect 418 244 426 261
rect 393 236 426 244
rect -42 215 116 217
rect -73 213 116 215
rect -73 205 246 213
rect -73 200 221 205
rect -73 199 -65 200
rect -98 191 -65 199
rect -42 197 221 200
rect -42 97 -27 197
rect 213 188 221 197
rect 238 188 246 205
rect 213 180 246 188
rect 101 160 134 168
rect 101 143 109 160
rect 126 143 134 160
rect 101 135 134 143
rect 101 97 116 135
rect 222 97 237 180
rect 393 97 408 236
rect 488 152 503 289
rect 621 260 654 267
rect 681 260 696 289
rect 802 267 817 289
rect 621 259 696 260
rect 621 242 629 259
rect 646 245 696 259
rect 646 242 654 245
rect 621 234 654 242
rect 681 213 696 245
rect 793 259 826 267
rect 793 242 801 259
rect 818 242 826 259
rect 793 234 826 242
rect 997 232 1012 289
rect 997 224 1030 232
rect 681 205 826 213
rect 681 197 801 205
rect 793 188 801 197
rect 818 188 826 205
rect 793 180 826 188
rect 997 207 1005 224
rect 1022 207 1030 224
rect 997 199 1030 207
rect 470 144 503 152
rect 470 127 478 144
rect 495 127 503 144
rect 470 119 503 127
rect 488 97 503 119
rect 681 160 714 168
rect 681 143 689 160
rect 706 143 714 160
rect 681 135 714 143
rect 681 97 696 135
rect 802 97 817 180
rect 997 97 1012 199
rect 1092 148 1107 289
rect 1074 140 1107 148
rect 1074 123 1082 140
rect 1099 123 1107 140
rect 1074 115 1107 123
rect 1092 97 1107 115
rect -42 40 -27 55
rect 101 40 116 55
rect 222 40 237 55
rect 393 40 408 55
rect 488 40 503 55
rect 681 40 696 55
rect 802 40 817 55
rect 997 40 1012 55
rect 1092 40 1107 55
<< polycont >>
rect -90 199 -73 216
rect 221 242 238 259
rect 401 244 418 261
rect 221 188 238 205
rect 109 143 126 160
rect 629 242 646 259
rect 801 242 818 259
rect 801 188 818 205
rect 1005 207 1022 224
rect 478 127 495 144
rect 689 143 706 160
rect 1082 123 1099 140
<< locali >>
rect -100 415 1165 423
rect -100 398 -70 415
rect -53 398 4 415
rect 21 398 73 415
rect 90 398 152 415
rect 169 398 225 415
rect 242 398 380 415
rect 397 398 459 415
rect 476 398 538 415
rect 555 398 653 415
rect 670 398 732 415
rect 749 398 805 415
rect 822 398 984 415
rect 1001 398 1063 415
rect 1080 398 1165 415
rect -100 390 1165 398
rect -80 334 -60 390
rect 436 334 456 390
rect 1040 334 1060 390
rect -86 326 -53 334
rect -86 309 -78 326
rect -61 309 -53 326
rect -86 301 -53 309
rect -17 326 16 334
rect -17 309 -9 326
rect 8 309 16 326
rect -17 301 16 309
rect 57 326 90 334
rect 57 309 65 326
rect 82 309 90 326
rect 57 301 90 309
rect 167 326 200 334
rect 167 309 175 326
rect 192 309 200 326
rect 167 301 200 309
rect 262 330 295 334
rect 350 330 383 334
rect 262 326 383 330
rect 262 309 270 326
rect 287 309 358 326
rect 375 309 383 326
rect 262 305 383 309
rect 262 301 295 305
rect 350 301 383 305
rect 433 326 466 334
rect 433 309 441 326
rect 458 309 466 326
rect 433 301 466 309
rect 508 326 670 334
rect 508 309 516 326
rect 533 309 645 326
rect 662 309 670 326
rect 508 301 670 309
rect 747 326 780 334
rect 747 309 755 326
rect 772 309 780 326
rect 747 301 780 309
rect 842 326 875 334
rect 842 309 850 326
rect 867 325 875 326
rect 946 326 979 334
rect 946 325 954 326
rect 867 309 954 325
rect 971 309 979 326
rect 842 305 979 309
rect 842 301 875 305
rect 946 301 979 305
rect 1037 326 1070 334
rect 1037 309 1045 326
rect 1062 309 1070 326
rect 1037 301 1070 309
rect 1112 326 1145 334
rect 1112 309 1120 326
rect 1137 309 1145 326
rect 1112 301 1145 309
rect -98 216 -65 224
rect -98 199 -90 216
rect -73 199 -65 216
rect -98 173 -65 199
rect -98 156 -90 173
rect -73 156 -65 173
rect -10 166 10 301
rect 60 261 80 301
rect 52 255 80 261
rect 52 238 57 255
rect 74 238 80 255
rect 52 233 80 238
rect -98 149 -65 156
rect -11 160 18 166
rect -11 143 -5 160
rect 12 143 18 160
rect -11 137 18 143
rect -10 94 10 137
rect 60 94 80 233
rect 101 160 134 168
rect 101 143 109 160
rect 126 143 134 160
rect 101 135 134 143
rect 172 155 192 301
rect 213 259 246 267
rect 213 242 221 259
rect 238 242 246 259
rect 213 234 246 242
rect 213 205 246 213
rect 213 188 221 205
rect 238 188 246 205
rect 213 180 246 188
rect 172 147 204 155
rect 172 130 180 147
rect 197 130 204 147
rect 172 124 204 130
rect 172 94 192 124
rect 267 94 287 301
rect 393 262 426 269
rect 521 262 541 301
rect 393 261 541 262
rect 393 244 401 261
rect 418 244 541 261
rect 393 242 541 244
rect 393 236 426 242
rect 470 144 503 152
rect 470 127 478 144
rect 495 127 503 144
rect 470 119 503 127
rect 521 94 541 242
rect 621 259 654 267
rect 621 242 629 259
rect 646 242 654 259
rect 621 234 654 242
rect 681 160 714 168
rect 681 143 689 160
rect 706 143 714 160
rect 681 135 714 143
rect 752 156 772 301
rect 793 259 826 267
rect 793 242 801 259
rect 818 242 826 259
rect 793 234 826 242
rect 793 205 826 213
rect 793 188 801 205
rect 818 188 826 205
rect 793 180 826 188
rect 752 148 784 156
rect 752 131 760 148
rect 777 131 784 148
rect 752 125 784 131
rect 752 94 772 125
rect 847 94 867 301
rect 939 225 1030 232
rect 1125 225 1145 301
rect 939 224 1145 225
rect 939 207 946 224
rect 963 207 1005 224
rect 1022 207 1145 224
rect 939 205 1145 207
rect 939 200 1030 205
rect 997 199 1030 200
rect 1074 140 1107 148
rect 1074 123 1082 140
rect 1099 123 1107 140
rect 1074 115 1107 123
rect 1125 94 1145 205
rect -86 86 -53 94
rect -86 69 -78 86
rect -61 69 -53 86
rect -86 61 -53 69
rect -17 86 16 94
rect -17 69 -9 86
rect 8 69 16 86
rect -17 61 16 69
rect 57 86 90 94
rect 57 69 65 86
rect 82 69 90 86
rect 57 61 90 69
rect 167 86 200 94
rect 167 69 175 86
rect 192 69 200 86
rect 167 61 200 69
rect 262 86 295 94
rect 262 69 270 86
rect 287 85 295 86
rect 345 85 378 93
rect 287 69 353 85
rect 262 68 353 69
rect 370 68 378 85
rect 262 65 378 68
rect 262 61 295 65
rect -80 14 -60 61
rect 345 60 378 65
rect 433 86 466 94
rect 433 69 441 86
rect 458 69 466 86
rect 433 61 466 69
rect 446 14 466 61
rect 508 86 670 94
rect 508 69 516 86
rect 533 69 645 86
rect 662 69 670 86
rect 508 60 670 69
rect 747 86 780 94
rect 747 69 755 86
rect 772 69 780 86
rect 747 61 780 69
rect 842 86 875 94
rect 842 69 850 86
rect 867 85 875 86
rect 949 86 982 94
rect 949 85 957 86
rect 867 69 957 85
rect 974 69 982 86
rect 842 65 982 69
rect 842 61 875 65
rect 949 61 982 65
rect 1037 86 1070 94
rect 1037 69 1045 86
rect 1062 69 1070 86
rect 1037 61 1070 69
rect 1112 86 1145 94
rect 1112 69 1120 86
rect 1137 69 1145 86
rect 1112 61 1145 69
rect 1050 14 1070 61
rect -106 6 1147 14
rect -106 -11 -91 6
rect -74 -11 -31 6
rect -14 -11 52 6
rect 69 -11 112 6
rect 129 -11 156 6
rect 173 -11 216 6
rect 233 -11 267 6
rect 284 -11 403 6
rect 420 -11 452 6
rect 469 -11 512 6
rect 529 -11 632 6
rect 649 -11 692 6
rect 709 -11 736 6
rect 753 -11 796 6
rect 813 -11 847 6
rect 864 -11 1007 6
rect 1024 -11 1056 6
rect 1073 -11 1116 6
rect 1133 -11 1147 6
rect -106 -19 1147 -11
<< viali >>
rect 4 398 21 415
rect 152 398 169 415
rect 380 398 397 415
rect 538 398 555 415
rect 732 398 749 415
rect 984 398 1001 415
rect -90 156 -73 173
rect 57 238 74 255
rect -5 143 12 160
rect 109 143 126 160
rect 221 242 238 259
rect 221 188 238 205
rect 180 130 197 147
rect 478 127 495 144
rect 629 242 646 259
rect 689 143 706 160
rect 801 242 818 259
rect 760 131 777 148
rect 946 207 963 224
rect 1082 123 1099 140
rect -31 -11 -14 6
rect 112 -11 129 6
rect 216 -11 233 6
rect 403 -11 420 6
rect 512 -11 529 6
rect 692 -11 709 6
rect 796 -11 813 6
rect 1007 -11 1024 6
rect 1116 -11 1133 6
<< metal1 >>
rect -106 415 1165 429
rect -106 398 4 415
rect 21 398 152 415
rect 169 398 380 415
rect 397 398 538 415
rect 555 398 732 415
rect 749 398 984 415
rect 1001 398 1165 415
rect -106 384 1165 398
rect 17 260 80 263
rect 17 234 21 260
rect 47 255 80 260
rect 213 259 246 267
rect 213 255 221 259
rect 47 238 57 255
rect 74 238 80 255
rect 47 234 80 238
rect 17 231 80 234
rect 105 242 221 255
rect 238 255 246 259
rect 621 259 654 267
rect 621 255 629 259
rect 238 242 629 255
rect 646 242 654 259
rect 793 259 826 267
rect 793 255 801 259
rect 105 235 654 242
rect -98 178 -30 181
rect -98 173 -59 178
rect -98 156 -90 173
rect -73 156 -59 173
rect -98 152 -59 156
rect -33 152 -30 178
rect 105 168 125 235
rect 213 234 246 235
rect 621 234 654 235
rect 685 242 801 255
rect 818 242 826 259
rect 685 235 826 242
rect 213 210 246 213
rect 685 210 705 235
rect 793 234 826 235
rect 213 205 705 210
rect 213 188 221 205
rect 238 188 705 205
rect 907 229 970 232
rect 907 203 910 229
rect 936 224 970 229
rect 936 207 946 224
rect 963 207 970 224
rect 936 203 970 207
rect 907 200 970 203
rect 213 185 705 188
rect 213 180 246 185
rect 685 168 705 185
rect -98 149 -30 152
rect -11 160 18 166
rect 101 160 134 168
rect -11 143 -5 160
rect 12 143 109 160
rect 126 143 134 160
rect 681 160 714 168
rect -11 140 134 143
rect -11 137 18 140
rect 101 135 134 140
rect 174 147 204 155
rect 174 130 180 147
rect 197 145 204 147
rect 470 145 503 152
rect 197 144 503 145
rect 197 130 478 144
rect 174 127 478 130
rect 495 127 503 144
rect 681 143 689 160
rect 706 143 714 160
rect 681 135 714 143
rect 754 148 784 156
rect 174 124 503 127
rect 754 131 760 148
rect 777 145 784 148
rect 1073 145 1107 148
rect 777 140 1107 145
rect 777 131 1082 140
rect 754 125 1082 131
rect 470 119 503 124
rect 1073 123 1082 125
rect 1099 123 1107 140
rect 1073 115 1107 123
rect -106 6 1165 20
rect -106 -11 -31 6
rect -14 -11 112 6
rect 129 -11 216 6
rect 233 -11 403 6
rect 420 -11 512 6
rect 529 -11 692 6
rect 709 -11 796 6
rect 813 -11 1007 6
rect 1024 -11 1116 6
rect 1133 -11 1165 6
rect -106 -25 1165 -11
<< via1 >>
rect 21 234 47 260
rect -59 152 -33 178
rect 910 203 936 229
<< metal2 >>
rect 17 260 51 263
rect 17 234 21 260
rect 47 234 51 260
rect 17 231 51 234
rect 907 229 939 232
rect 907 203 910 229
rect 936 203 939 229
rect 907 200 939 203
rect -61 178 -30 181
rect -61 152 -59 178
rect -33 152 -30 178
rect -61 149 -30 152
<< labels >>
flabel metal2 s 21 234 47 260 0 FreeSans 400 0 0 0 D
port 2 nsew
flabel locali s 183 134 191 141 0 FreeSans 200 0 0 0 net1
flabel locali s 273 160 281 168 0 FreeSans 200 0 0 0 net2
flabel metal1 s 486 396 525 416 0 FreeSans 400 0 0 0 vdd
port 0 nsew
flabel metal1 s 433 -19 568 14 0 FreeSans 400 0 0 0 gnd
port 1 nsew
flabel locali s 529 128 537 136 0 FreeSans 200 0 0 0 net3
flabel locali s 765 134 773 141 0 FreeSans 200 0 0 0 net4
flabel locali s 852 310 862 322 0 FreeSans 200 0 0 0 net5
flabel metal2 s 910 203 936 229 0 FreeSans 400 0 0 0 Q
port 9 nsew
flabel metal2 s -59 152 -33 178 0 FreeSans 240 0 0 0 clk
port 10 nsew
flabel locali s 111 144 122 157 0 FreeSans 240 0 0 0 clkb
<< properties >>
string FIXED_BBOX -106 -3 1165 406
<< end >>
