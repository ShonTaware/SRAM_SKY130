magic
tech sky130A
timestamp 1615985747
<< nwell >>
rect -3 425 483 677
rect -3 424 81 425
<< nmos >>
rect 60 290 75 332
rect 193 290 208 332
rect 328 325 343 367
rect 423 303 465 318
<< pmos >>
rect 60 445 75 571
rect 193 445 208 571
rect 328 445 343 500
<< ndiff >>
rect 283 358 328 367
rect 283 341 296 358
rect 313 341 328 358
rect 15 322 60 332
rect 15 305 28 322
rect 45 305 60 322
rect 15 290 60 305
rect 75 322 120 332
rect 75 305 90 322
rect 107 305 120 322
rect 75 290 120 305
rect 148 322 193 332
rect 148 305 161 322
rect 178 305 193 322
rect 148 290 193 305
rect 208 322 253 332
rect 283 325 328 341
rect 343 359 388 367
rect 343 342 358 359
rect 375 342 388 359
rect 343 325 388 342
rect 208 305 223 322
rect 240 305 253 322
rect 423 350 465 363
rect 423 333 438 350
rect 455 333 465 350
rect 423 318 465 333
rect 208 290 253 305
rect 423 288 465 303
rect 423 271 438 288
rect 455 271 465 288
rect 423 258 465 271
<< pdiff >>
rect 15 557 60 571
rect 15 540 29 557
rect 46 540 60 557
rect 15 484 60 540
rect 15 467 29 484
rect 46 467 60 484
rect 15 445 60 467
rect 75 551 121 571
rect 75 534 90 551
rect 107 534 121 551
rect 75 484 121 534
rect 75 467 90 484
rect 107 467 121 484
rect 75 445 121 467
rect 148 557 193 571
rect 148 540 162 557
rect 179 540 193 557
rect 148 484 193 540
rect 148 467 162 484
rect 179 467 193 484
rect 148 445 193 467
rect 208 551 254 571
rect 208 534 223 551
rect 240 534 254 551
rect 208 484 254 534
rect 208 467 223 484
rect 240 467 254 484
rect 208 445 254 467
rect 283 484 328 500
rect 283 467 297 484
rect 314 467 328 484
rect 283 445 328 467
rect 343 484 389 500
rect 343 467 358 484
rect 375 467 389 484
rect 343 445 389 467
<< ndiffc >>
rect 296 341 313 358
rect 28 305 45 322
rect 90 305 107 322
rect 161 305 178 322
rect 358 342 375 359
rect 223 305 240 322
rect 438 333 455 350
rect 438 271 455 288
<< pdiffc >>
rect 29 540 46 557
rect 29 467 46 484
rect 90 534 107 551
rect 90 467 107 484
rect 162 540 179 557
rect 162 467 179 484
rect 223 534 240 551
rect 223 467 240 484
rect 297 467 314 484
rect 358 467 375 484
<< psubdiff >>
rect 48 232 89 244
rect 48 215 60 232
rect 77 215 89 232
rect 48 203 89 215
rect 181 232 222 244
rect 181 215 193 232
rect 210 215 222 232
rect 181 203 222 215
rect 316 232 357 244
rect 316 215 328 232
rect 345 215 357 232
rect 316 203 357 215
<< nsubdiff >>
rect 72 634 125 652
rect 72 617 90 634
rect 107 617 125 634
rect 72 599 125 617
rect 205 634 258 652
rect 205 617 223 634
rect 240 617 258 634
rect 205 599 258 617
rect 340 634 393 652
rect 340 617 358 634
rect 375 617 393 634
rect 340 599 393 617
<< psubdiffcont >>
rect 60 215 77 232
rect 193 215 210 232
rect 328 215 345 232
<< nsubdiffcont >>
rect 90 617 107 634
rect 223 617 240 634
rect 358 617 375 634
<< poly >>
rect 60 571 75 585
rect 193 571 208 585
rect 320 570 353 578
rect 320 553 328 570
rect 345 553 353 570
rect 320 545 353 553
rect 328 500 343 545
rect 5 389 38 397
rect 5 372 13 389
rect 30 385 38 389
rect 60 385 75 445
rect 30 372 75 385
rect 5 370 75 372
rect 5 364 38 370
rect 60 332 75 370
rect 139 389 172 397
rect 139 372 147 389
rect 164 385 172 389
rect 193 385 208 445
rect 328 433 343 445
rect 328 418 413 433
rect 164 372 208 385
rect 139 370 208 372
rect 139 364 172 370
rect 193 332 208 370
rect 328 367 343 380
rect 328 313 343 325
rect 397 318 413 418
rect 319 305 352 313
rect 60 277 75 290
rect 193 277 208 290
rect 319 288 327 305
rect 344 288 352 305
rect 397 303 423 318
rect 465 303 483 318
rect 319 280 352 288
<< polycont >>
rect 328 553 345 570
rect 13 372 30 389
rect 147 372 164 389
rect 327 288 344 305
<< locali >>
rect -3 635 483 642
rect -3 618 38 635
rect 55 634 171 635
rect 55 618 90 634
rect -3 617 90 618
rect 107 618 171 634
rect 188 634 251 635
rect 188 618 223 634
rect 107 617 223 618
rect 240 618 251 634
rect 268 618 306 635
rect 323 634 416 635
rect 323 618 358 634
rect 240 617 358 618
rect 375 618 416 634
rect 433 618 483 635
rect 375 617 483 618
rect -3 609 483 617
rect 19 557 55 609
rect 19 540 29 557
rect 46 540 55 557
rect 19 484 55 540
rect 19 467 29 484
rect 46 467 55 484
rect 19 445 55 467
rect 82 551 115 561
rect 82 534 90 551
rect 107 534 115 551
rect 82 484 115 534
rect 82 467 90 484
rect 107 467 115 484
rect 5 390 38 397
rect 4 389 38 390
rect 4 372 13 389
rect 30 372 38 389
rect 4 370 38 372
rect 5 364 38 370
rect 82 390 115 467
rect 152 557 188 609
rect 320 570 353 578
rect 152 540 162 557
rect 179 540 188 557
rect 152 484 188 540
rect 152 467 162 484
rect 179 467 188 484
rect 152 445 188 467
rect 215 551 248 561
rect 215 534 223 551
rect 240 534 248 551
rect 320 553 328 570
rect 345 553 353 570
rect 320 545 353 553
rect 215 484 248 534
rect 215 467 223 484
rect 240 467 248 484
rect 139 390 172 397
rect 82 389 172 390
rect 82 372 147 389
rect 164 372 172 389
rect 82 370 172 372
rect 20 322 53 330
rect 20 305 28 322
rect 45 305 53 322
rect 20 240 53 305
rect 82 322 115 370
rect 139 364 172 370
rect 215 360 248 467
rect 287 484 323 500
rect 287 467 297 484
rect 314 467 323 484
rect 287 445 323 467
rect 350 484 383 500
rect 350 467 358 484
rect 375 467 383 484
rect 297 367 317 445
rect 288 360 321 367
rect 215 358 321 360
rect 215 341 296 358
rect 313 341 321 358
rect 215 340 321 341
rect 82 305 90 322
rect 107 305 115 322
rect 82 297 115 305
rect 153 322 186 330
rect 153 305 161 322
rect 178 305 186 322
rect 153 240 186 305
rect 215 322 248 340
rect 288 331 321 340
rect 350 359 383 467
rect 350 342 358 359
rect 375 355 383 359
rect 423 355 463 358
rect 375 350 463 355
rect 375 342 438 350
rect 350 335 438 342
rect 350 331 383 335
rect 423 333 438 335
rect 455 333 463 350
rect 423 325 463 333
rect 215 305 223 322
rect 240 305 248 322
rect 215 297 248 305
rect 319 305 352 313
rect 319 288 327 305
rect 344 288 352 305
rect 319 280 352 288
rect 430 288 465 296
rect 430 271 438 288
rect 455 271 465 288
rect 430 263 465 271
rect 434 240 458 263
rect -3 232 483 240
rect -3 215 60 232
rect 77 215 193 232
rect 210 215 253 232
rect 270 215 328 232
rect 345 215 403 232
rect 420 215 483 232
rect -3 207 483 215
<< viali >>
rect 38 618 55 635
rect 171 618 188 635
rect 251 618 268 635
rect 306 618 323 635
rect 416 618 433 635
rect 253 215 270 232
rect 403 215 420 232
<< metal1 >>
rect -3 635 483 648
rect -3 618 38 635
rect 55 618 171 635
rect 188 618 251 635
rect 268 618 306 635
rect 323 618 416 635
rect 433 618 483 635
rect -3 598 483 618
rect -3 232 483 250
rect -3 215 253 232
rect 270 215 403 232
rect 420 215 483 232
rect -3 200 483 215
<< labels >>
flabel metal1 s 156 211 207 234 7 FreeSans 200 0 0 0 gnd
port 11 w
flabel locali s 15 373 26 386 7 FreeSans 400 0 0 0 in
port 1 w
flabel locali s 232 346 259 356 0 FreeSans 200 0 0 0 net2
flabel locali s 144 375 175 385 7 FreeSans 200 0 0 0 net1
flabel locali s 359 385 369 395 0 FreeSans 200 0 0 0 out
port 13 nsew
flabel locali s 325 284 347 306 7 FreeSans 400 0 0 0 en
port 4 w
flabel metal1 s 156 602 279 645 7 FreeSans 200 0 0 0 vdd
port 12 w
flabel locali s 325 549 347 571 7 FreeSans 400 0 0 0 enb
port 5 w
<< properties >>
string FIXED_BBOX -3 223 483 625
<< end >>
