

.lib "./sky130.lib.spice" ff

