Sense Amplifier

.lib "./libs/models/sky130.lib.spice" tt

XM1 net1 blb net2 gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.21
XM3 out bl net2 gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.21

XM2 net1 net1 vdd vdd sky130_fd_pr__pfet_01v8 w=0.42 l=0.21
XM4 out net1 vdd vdd sky130_fd_pr__pfet_01v8 w=0.84 l=0.21

XM5 net2 rd_en gnd gnd sky130_fd_pr__nfet_01v8 w=1.26 l=0.21

XM6 dout out gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.21
XM7 dout out vdd vdd sky130_fd_pr__pfet_01v8 w=0.42 l=0.21

V1 vdd gnd dc 1.8v
V2 blb 0 pulse 1.8 0 0 60ps 60ps 1ns 2ns
V3 bl 0 pulse 0 1.8 0 60ps 60ps 1ns 2ns
V4 rd_en 0 pulse 0 1.8 0 60ps 60ps 5ns 10ns

.tran 0.1p 20n
.control
run
plot V(rd_en)+6 V(bl)+4 V(blb)+2 V(dout) 
.endc
.end


